magic
tech sky130A
magscale 1 2
timestamp 1713067979
<< pwell >>
rect -683 -1010 683 1010
<< nmos >>
rect -487 -800 -287 800
rect -229 -800 -29 800
rect 29 -800 229 800
rect 287 -800 487 800
<< ndiff >>
rect -545 788 -487 800
rect -545 -788 -533 788
rect -499 -788 -487 788
rect -545 -800 -487 -788
rect -287 788 -229 800
rect -287 -788 -275 788
rect -241 -788 -229 788
rect -287 -800 -229 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 229 788 287 800
rect 229 -788 241 788
rect 275 -788 287 788
rect 229 -800 287 -788
rect 487 788 545 800
rect 487 -788 499 788
rect 533 -788 545 788
rect 487 -800 545 -788
<< ndiffc >>
rect -533 -788 -499 788
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect 499 -788 533 788
<< psubdiff >>
rect -647 940 647 974
rect -647 878 -613 940
rect 613 878 647 940
rect -647 -940 -613 -878
rect 613 -940 647 -878
rect -647 -974 -551 -940
rect 551 -974 647 -940
<< psubdiffcont >>
rect -647 -878 -613 878
rect 613 -878 647 878
rect -551 -974 551 -940
<< poly >>
rect -487 872 -287 888
rect -487 838 -471 872
rect -303 838 -287 872
rect -487 800 -287 838
rect -229 872 -29 888
rect -229 838 -213 872
rect -45 838 -29 872
rect -229 800 -29 838
rect 29 872 229 888
rect 29 838 45 872
rect 213 838 229 872
rect 29 800 229 838
rect 287 872 487 888
rect 287 838 303 872
rect 471 838 487 872
rect 287 800 487 838
rect -487 -838 -287 -800
rect -487 -872 -471 -838
rect -303 -872 -287 -838
rect -487 -888 -287 -872
rect -229 -838 -29 -800
rect -229 -872 -213 -838
rect -45 -872 -29 -838
rect -229 -888 -29 -872
rect 29 -838 229 -800
rect 29 -872 45 -838
rect 213 -872 229 -838
rect 29 -888 229 -872
rect 287 -838 487 -800
rect 287 -872 303 -838
rect 471 -872 487 -838
rect 287 -888 487 -872
<< polycont >>
rect -471 838 -303 872
rect -213 838 -45 872
rect 45 838 213 872
rect 303 838 471 872
rect -471 -872 -303 -838
rect -213 -872 -45 -838
rect 45 -872 213 -838
rect 303 -872 471 -838
<< locali >>
rect -647 878 -613 974
rect 613 878 647 974
rect -487 838 -471 872
rect -303 838 -287 872
rect -229 838 -213 872
rect -45 838 -29 872
rect 29 838 45 872
rect 213 838 229 872
rect 287 838 303 872
rect 471 838 487 872
rect -533 788 -499 804
rect -533 -804 -499 -788
rect -275 788 -241 804
rect -275 -804 -241 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 241 788 275 804
rect 241 -804 275 -788
rect 499 788 533 804
rect 499 -804 533 -788
rect -487 -872 -471 -838
rect -303 -872 -287 -838
rect -229 -872 -213 -838
rect -45 -872 -29 -838
rect 29 -872 45 -838
rect 213 -872 229 -838
rect 287 -872 303 -838
rect 471 -872 487 -838
rect -647 -974 -551 -940
rect 551 -974 647 -940
<< viali >>
rect -613 940 613 974
rect -471 838 -303 872
rect -213 838 -45 872
rect 45 838 213 872
rect 303 838 471 872
rect -647 -878 -613 -188
rect -533 141 -499 771
rect -275 -771 -241 -141
rect -17 141 17 771
rect 241 -771 275 -141
rect 499 141 533 771
rect -471 -872 -303 -838
rect -213 -872 -45 -838
rect 45 -872 213 -838
rect 303 -872 471 -838
rect -647 -940 -613 -878
rect 613 -878 647 -188
rect 613 -940 647 -878
<< metal1 >>
rect -625 974 625 980
rect -625 940 -613 974
rect 613 940 625 974
rect -625 934 625 940
rect -483 872 -291 878
rect -483 838 -471 872
rect -303 838 -291 872
rect -483 832 -291 838
rect -225 872 -33 878
rect -225 838 -213 872
rect -45 838 -33 872
rect -225 832 -33 838
rect 33 872 225 878
rect 33 838 45 872
rect 213 838 225 872
rect 33 832 225 838
rect 291 872 483 878
rect 291 838 303 872
rect 471 838 483 872
rect 291 832 483 838
rect -539 771 -493 783
rect -539 141 -533 771
rect -499 141 -493 771
rect -539 129 -493 141
rect -23 771 23 783
rect -23 141 -17 771
rect 17 141 23 771
rect -23 129 23 141
rect 493 771 539 783
rect 493 141 499 771
rect 533 141 539 771
rect 493 129 539 141
rect -281 -141 -235 -129
rect -653 -188 -607 -176
rect -653 -940 -647 -188
rect -613 -940 -607 -188
rect -281 -771 -275 -141
rect -241 -771 -235 -141
rect -281 -783 -235 -771
rect 235 -141 281 -129
rect 235 -771 241 -141
rect 275 -771 281 -141
rect 235 -783 281 -771
rect 607 -188 653 -176
rect -483 -838 -291 -832
rect -483 -872 -471 -838
rect -303 -872 -291 -838
rect -483 -878 -291 -872
rect -225 -838 -33 -832
rect -225 -872 -213 -838
rect -45 -872 -33 -838
rect -225 -878 -33 -872
rect 33 -838 225 -832
rect 33 -872 45 -838
rect 213 -872 225 -838
rect 33 -878 225 -872
rect 291 -838 483 -832
rect 291 -872 303 -838
rect 471 -872 483 -838
rect 291 -878 483 -872
rect -653 -952 -607 -940
rect 607 -940 613 -188
rect 647 -940 653 -188
rect 607 -952 653 -940
<< properties >>
string FIXED_BBOX -630 -957 630 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
