magic
tech sky130A
magscale 1 2
timestamp 1713485453
<< metal1 >>
rect 29638 4278 29938 4308
rect 29632 3978 29638 4278
rect 29938 3978 29944 4278
rect 29638 3664 29938 3978
rect 28886 3364 29938 3664
rect 29974 3196 30094 3202
rect 29630 3184 29974 3196
rect 29046 3076 29974 3184
rect 31354 3184 31494 3190
rect 30094 3076 31354 3184
rect 29046 3044 31354 3076
rect 31354 3038 31494 3044
rect 10908 1740 11976 2138
rect 29086 1764 29598 1864
rect 10908 1451 11334 1740
rect 11623 1451 11976 1740
rect 10908 1264 11976 1451
rect 11334 1203 11623 1264
rect 11334 1150 28017 1203
rect 29032 1150 29152 1204
rect 11334 914 29152 1150
rect 27722 912 29152 914
rect 29499 806 29598 1764
rect 29493 707 29499 806
rect 29598 707 29604 806
<< via1 >>
rect 29638 3978 29938 4278
rect 29974 3076 30094 3196
rect 31354 3044 31494 3184
rect 11334 1451 11623 1740
rect 29499 707 29598 806
<< metal2 >>
rect 29638 4278 29938 4284
rect 29629 3978 29638 4278
rect 29938 3978 29947 4278
rect 29638 3972 29938 3978
rect 29968 3076 29974 3196
rect 30094 3193 31432 3196
rect 30094 3191 31494 3193
rect 30094 3081 31317 3191
rect 31427 3184 31494 3191
rect 30094 3076 31354 3081
rect 31348 3044 31354 3076
rect 31494 3044 31500 3184
rect 31354 3035 31494 3044
rect 10908 1740 11976 2138
rect 10908 1451 11334 1740
rect 11623 1451 11976 1740
rect 10908 1264 11976 1451
rect 29499 806 29598 812
rect 29490 707 29499 806
rect 29598 707 29607 806
rect 29499 701 29598 707
<< via2 >>
rect 29638 3978 29938 4278
rect 31317 3184 31427 3191
rect 31317 3081 31354 3184
rect 31354 3044 31494 3184
rect 11334 1451 11623 1740
rect 29499 707 29598 806
<< metal3 >>
rect 29633 4278 29943 4283
rect 26862 4277 29638 4278
rect 1754 3980 1760 4277
rect 2057 3980 29638 4277
rect 26862 3978 29638 3980
rect 29938 3978 29943 4278
rect 29633 3973 29943 3978
rect 31313 3196 31431 3201
rect 31312 3195 31432 3196
rect 31312 3077 31313 3195
rect 31431 3189 31432 3195
rect 31431 3184 31499 3189
rect 31312 3076 31354 3077
rect 31313 3071 31354 3076
rect 31349 3044 31354 3071
rect 31494 3044 31499 3184
rect 31349 3039 31499 3044
rect 10908 2012 11976 2138
rect 10716 1740 11976 2012
rect 9798 1451 9804 1740
rect 10093 1451 11334 1740
rect 11623 1451 11976 1740
rect 10716 1264 11976 1451
rect 31354 1338 31494 3039
rect 10716 1242 11920 1264
rect 29488 702 29494 811
rect 29593 806 29603 811
rect 29598 707 29603 806
rect 29593 702 29603 707
<< via3 >>
rect 1760 3980 2057 4277
rect 31313 3191 31431 3195
rect 31313 3081 31317 3191
rect 31317 3184 31427 3191
rect 31427 3184 31431 3191
rect 31317 3081 31431 3184
rect 31313 3077 31354 3081
rect 31354 3077 31431 3081
rect 9804 1451 10093 1740
rect 29494 806 29593 811
rect 29494 707 29499 806
rect 29499 707 29593 806
rect 29494 702 29593 707
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 4277 500 44152
rect 1759 4277 2058 4278
rect 180 3980 1760 4277
rect 2057 3980 2058 4277
rect 200 1000 500 3980
rect 1759 3979 2058 3980
rect 9800 1740 10100 44152
rect 9800 1451 9804 1740
rect 10093 1451 10100 1740
rect 9800 1000 10100 1451
rect 31312 3195 31432 3196
rect 31312 3077 31313 3195
rect 31431 3077 31432 3195
rect 29493 811 29594 812
rect 29493 806 29494 811
rect 26911 707 29494 806
rect 26911 200 27010 707
rect 29493 702 29494 707
rect 29593 702 29594 811
rect 29493 701 29594 702
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 3077
use idac1  idac1_0
timestamp 1713485344
transform 0 -1 18130 1 0 15144
box 0 -2600 9600 2600
use opamp1  opamp1_0
timestamp 1713144495
transform 1 0 22231 0 1 7854
box 1445 -1430 5650 2100
use vbias1  vbias1_0
timestamp 1713046980
transform 1 0 21530 0 1 7912
box -400 -640 1060 1968
use vbias1  vbias1_1
timestamp 1713046980
transform 1 0 28126 0 1 1724
box -400 -640 1060 1968
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
