magic
tech sky130A
magscale 1 2
timestamp 1725240473
<< metal1 >>
rect 0 2600 4160 2620
rect 0 2480 840 2600
rect 960 2480 4160 2600
rect 0 2440 4160 2480
rect 70 2040 80 2100
rect 140 2040 150 2100
rect 1270 2040 1280 2100
rect 1340 2040 1350 2100
rect 2550 2000 2560 2060
rect 2620 2000 2630 2060
rect 3030 2000 3040 2060
rect 3100 2000 3110 2060
rect 3510 2000 3520 2060
rect 3580 2000 3590 2060
rect 670 1900 680 1960
rect 740 1900 750 1960
rect 1870 1900 1880 1960
rect 1940 1900 1950 1960
rect 2730 1800 2740 1860
rect 2800 1800 2810 1860
rect 3210 1800 3220 1860
rect 3280 1800 3290 1860
rect 3690 1800 3700 1860
rect 3760 1800 3770 1860
rect -200 1340 3400 1460
rect 3520 1340 3820 1460
rect -200 1320 3820 1340
rect -200 100 -60 1320
rect 3980 1240 4160 2440
rect 0 1220 4160 1240
rect 0 1100 860 1220
rect 980 1100 4160 1220
rect 0 1080 4160 1100
rect 70 680 80 740
rect 140 680 150 740
rect 1270 680 1280 740
rect 1340 680 1350 740
rect 2470 680 2480 740
rect 2540 680 2550 740
rect 670 540 680 600
rect 740 540 750 600
rect 1870 540 1880 600
rect 1940 540 1950 600
rect 2860 540 3140 600
rect 3320 540 3610 600
rect 3740 420 3750 500
rect 3830 420 3840 500
rect 3370 100 3380 140
rect -200 20 3380 100
rect 3500 100 3510 140
rect 3500 20 3980 100
rect -200 0 3980 20
<< via1 >>
rect 840 2480 960 2600
rect 80 2040 140 2100
rect 1280 2040 1340 2100
rect 2560 2000 2620 2060
rect 3040 2000 3100 2060
rect 3520 2000 3580 2060
rect 680 1900 740 1960
rect 1880 1900 1940 1960
rect 2740 1800 2800 1860
rect 3220 1800 3280 1860
rect 3700 1800 3760 1860
rect 3400 1340 3520 1460
rect 860 1100 980 1220
rect 80 680 140 740
rect 1280 680 1340 740
rect 2480 680 2540 740
rect 680 540 740 600
rect 1880 540 1940 600
rect 3750 420 3830 500
rect 3380 20 3500 140
<< metal2 >>
rect 840 2600 960 2610
rect 840 2470 960 2480
rect 80 2100 880 2140
rect 140 2080 880 2100
rect 80 2030 140 2040
rect 440 1980 520 1990
rect 680 1960 740 1970
rect 520 1900 680 1960
rect 820 1920 880 2080
rect 1280 2100 2080 2140
rect 1340 2080 2080 2100
rect 1280 2030 1340 2040
rect 1680 1960 1740 1970
rect 1880 1960 1940 1970
rect 440 1890 520 1900
rect 680 1890 740 1900
rect 1740 1900 1880 1960
rect 2020 1920 2080 2080
rect 2560 2060 2620 2070
rect 3040 2060 3100 2070
rect 3520 2060 3580 2070
rect 2620 2000 3040 2060
rect 3100 2000 3520 2060
rect 3580 2000 3960 2060
rect 2560 1980 3960 2000
rect 1680 1890 1740 1900
rect 1880 1890 1940 1900
rect 20 1860 80 1870
rect 1300 1860 1360 1870
rect 2740 1860 2800 1870
rect 3220 1860 3280 1870
rect 3700 1860 3760 1870
rect 20 1790 80 1800
rect 940 1560 1020 1820
rect 1300 1790 1360 1800
rect 1800 1800 2740 1860
rect 2800 1800 3220 1860
rect 3280 1800 3700 1860
rect 3760 1800 3780 1860
rect 1800 1780 3780 1800
rect 1800 1560 1880 1780
rect 940 1480 1880 1560
rect 3400 1460 3520 1470
rect 3360 1340 3400 1460
rect 3520 1340 3560 1460
rect 860 1220 980 1230
rect 860 1090 980 1100
rect 80 740 880 780
rect 140 720 880 740
rect 80 670 140 680
rect 20 620 80 630
rect 80 560 260 620
rect 680 600 740 610
rect 20 550 80 560
rect 480 540 680 600
rect 820 560 880 720
rect 1280 740 2080 780
rect 2480 740 2540 750
rect 1340 720 2080 740
rect 1280 670 1340 680
rect 1320 620 1380 630
rect 680 530 740 540
rect 460 460 520 470
rect 520 400 680 460
rect 460 390 520 400
rect 1080 220 1140 580
rect 1380 560 1480 620
rect 1880 600 1940 610
rect 1320 550 1380 560
rect 1680 540 1880 600
rect 2020 560 2080 720
rect 2300 680 2480 740
rect 2300 540 2360 680
rect 2480 670 2540 680
rect 1880 530 1940 540
rect 1700 480 1880 500
rect 1760 420 1880 480
rect 1700 410 1760 420
rect 2400 220 2460 500
rect 1080 160 2460 220
rect 3360 140 3560 1340
rect 3880 520 3960 1980
rect 3750 500 3960 520
rect 3830 420 3960 500
rect 3750 410 3830 420
rect 3360 20 3380 140
rect 3500 20 3560 140
rect 3360 0 3560 20
<< via2 >>
rect 840 2480 960 2600
rect 440 1900 520 1980
rect 1680 1900 1740 1960
rect 20 1800 80 1860
rect 1300 1800 1360 1860
rect 860 1100 980 1220
rect 20 560 80 620
rect 460 400 520 460
rect 1320 560 1380 620
rect 1700 420 1760 480
<< metal3 >>
rect 820 2600 1020 2620
rect 820 2480 840 2600
rect 960 2480 1020 2600
rect 430 1980 530 1985
rect 20 1865 100 1920
rect 430 1900 440 1980
rect 520 1900 530 1980
rect 430 1895 530 1900
rect 10 1860 100 1865
rect 10 1800 20 1860
rect 80 1800 100 1860
rect 10 1795 100 1800
rect 20 625 100 1795
rect 10 620 100 625
rect 10 560 20 620
rect 80 560 100 620
rect 10 555 90 560
rect 440 465 520 1895
rect 820 1220 1020 2480
rect 1680 1965 1760 2000
rect 1670 1960 1760 1965
rect 1670 1900 1680 1960
rect 1740 1900 1760 1960
rect 1670 1895 1760 1900
rect 1290 1860 1370 1865
rect 1290 1800 1300 1860
rect 1360 1800 1380 1860
rect 1290 1795 1380 1800
rect 820 1100 860 1220
rect 980 1100 1020 1220
rect 820 1080 1020 1100
rect 1300 625 1380 1795
rect 1300 620 1390 625
rect 1300 560 1320 620
rect 1380 560 1390 620
rect 1300 555 1390 560
rect 1300 540 1380 555
rect 1680 485 1760 1895
rect 1680 480 1770 485
rect 440 460 530 465
rect 440 400 460 460
rect 520 400 530 460
rect 1680 420 1700 480
rect 1760 420 1770 480
rect 1680 415 1770 420
rect 1680 400 1760 415
rect 440 395 530 400
rect 440 380 520 395
use pll_inv1  pll_inv1_0
timestamp 1723400719
transform 1 0 3110 0 1 60
box -110 -60 390 1120
use pll_inv1  pll_inv1_1
timestamp 1723400719
transform 1 0 3050 0 1 1420
box -110 -60 390 1120
use pll_inv1  pll_inv1_2
timestamp 1723400719
transform 1 0 3590 0 1 60
box -110 -60 390 1120
use pll_inv1  pll_inv1_3
timestamp 1723400719
transform 1 0 2570 0 1 1420
box -110 -60 390 1120
use pll_inv1  pll_inv1_4
timestamp 1723400719
transform 1 0 3530 0 1 1420
box -110 -60 390 1120
use pll_nand  pll_nand_0
timestamp 1723401136
transform 1 0 2510 0 1 60
box -110 -60 550 1120
use pll_nor  pll_nor_0
timestamp 1723400899
transform 1 0 710 0 1 1420
box -110 -60 550 1120
use pll_nor  pll_nor_1
timestamp 1723400899
transform 1 0 110 0 1 1420
box -110 -60 550 1120
use pll_nor  pll_nor_2
timestamp 1723400899
transform 1 0 1910 0 1 1420
box -110 -60 550 1120
use pll_nor  pll_nor_3
timestamp 1723400899
transform 1 0 1310 0 1 1420
box -110 -60 550 1120
use pll_nor  pll_nor_4
timestamp 1723400899
transform 1 0 1310 0 1 60
box -110 -60 550 1120
use pll_nor  pll_nor_5
timestamp 1723400899
transform 1 0 1910 0 1 60
box -110 -60 550 1120
use pll_nor  pll_nor_6
timestamp 1723400899
transform 1 0 710 0 1 60
box -110 -60 550 1120
use pll_nor  pll_nor_7
timestamp 1723400899
transform 1 0 110 0 1 60
box -110 -60 550 1120
<< labels >>
flabel metal2 20 440 80 500 0 FreeSans 960 0 0 0 A
port 0 nsew
flabel metal2 1210 440 1270 500 0 FreeSans 960 0 0 0 B
port 1 nsew
flabel metal2 2400 160 2460 220 0 FreeSans 640 0 0 0 QA
port 2 nsew
flabel metal2 2300 680 2360 740 0 FreeSans 640 0 0 0 QB
port 3 nsew
flabel metal2 2920 1780 3000 1860 0 FreeSans 640 0 0 0 R
port 4 nsew
flabel metal2 620 540 680 600 0 FreeSans 640 0 0 0 QAB
flabel metal2 1820 540 1880 600 0 FreeSans 640 0 0 0 QBB
flabel metal2 1090 1900 1150 1920 0 FreeSans 640 0 0 0 RAB
flabel metal2 2290 1900 2350 1920 0 FreeSans 640 0 0 0 RBB
flabel metal1 0 0 100 100 0 FreeSans 1280 0 0 0 VSS
port 5 nsew
flabel metal1 0 2440 100 2540 0 FreeSans 1280 0 0 0 VDD
port 6 nsew
flabel metal2 2150 380 2210 440 0 FreeSans 640 0 0 0 RB
flabel metal2 950 380 1010 440 0 FreeSans 640 0 0 0 RA
<< end >>
