magic
tech sky130A
magscale 1 2
timestamp 1725372531
<< nwell >>
rect -1681 -615 1681 615
<< mvpmos >>
rect -1423 118 -1223 318
rect -1045 118 -845 318
rect -667 118 -467 318
rect -289 118 -89 318
rect 89 118 289 318
rect 467 118 667 318
rect 845 118 1045 318
rect 1223 118 1423 318
rect -1423 -318 -1223 -118
rect -1045 -318 -845 -118
rect -667 -318 -467 -118
rect -289 -318 -89 -118
rect 89 -318 289 -118
rect 467 -318 667 -118
rect 845 -318 1045 -118
rect 1223 -318 1423 -118
<< mvpdiff >>
rect -1481 306 -1423 318
rect -1481 130 -1469 306
rect -1435 130 -1423 306
rect -1481 118 -1423 130
rect -1223 306 -1165 318
rect -1223 130 -1211 306
rect -1177 130 -1165 306
rect -1223 118 -1165 130
rect -1103 306 -1045 318
rect -1103 130 -1091 306
rect -1057 130 -1045 306
rect -1103 118 -1045 130
rect -845 306 -787 318
rect -845 130 -833 306
rect -799 130 -787 306
rect -845 118 -787 130
rect -725 306 -667 318
rect -725 130 -713 306
rect -679 130 -667 306
rect -725 118 -667 130
rect -467 306 -409 318
rect -467 130 -455 306
rect -421 130 -409 306
rect -467 118 -409 130
rect -347 306 -289 318
rect -347 130 -335 306
rect -301 130 -289 306
rect -347 118 -289 130
rect -89 306 -31 318
rect -89 130 -77 306
rect -43 130 -31 306
rect -89 118 -31 130
rect 31 306 89 318
rect 31 130 43 306
rect 77 130 89 306
rect 31 118 89 130
rect 289 306 347 318
rect 289 130 301 306
rect 335 130 347 306
rect 289 118 347 130
rect 409 306 467 318
rect 409 130 421 306
rect 455 130 467 306
rect 409 118 467 130
rect 667 306 725 318
rect 667 130 679 306
rect 713 130 725 306
rect 667 118 725 130
rect 787 306 845 318
rect 787 130 799 306
rect 833 130 845 306
rect 787 118 845 130
rect 1045 306 1103 318
rect 1045 130 1057 306
rect 1091 130 1103 306
rect 1045 118 1103 130
rect 1165 306 1223 318
rect 1165 130 1177 306
rect 1211 130 1223 306
rect 1165 118 1223 130
rect 1423 306 1481 318
rect 1423 130 1435 306
rect 1469 130 1481 306
rect 1423 118 1481 130
rect -1481 -130 -1423 -118
rect -1481 -306 -1469 -130
rect -1435 -306 -1423 -130
rect -1481 -318 -1423 -306
rect -1223 -130 -1165 -118
rect -1223 -306 -1211 -130
rect -1177 -306 -1165 -130
rect -1223 -318 -1165 -306
rect -1103 -130 -1045 -118
rect -1103 -306 -1091 -130
rect -1057 -306 -1045 -130
rect -1103 -318 -1045 -306
rect -845 -130 -787 -118
rect -845 -306 -833 -130
rect -799 -306 -787 -130
rect -845 -318 -787 -306
rect -725 -130 -667 -118
rect -725 -306 -713 -130
rect -679 -306 -667 -130
rect -725 -318 -667 -306
rect -467 -130 -409 -118
rect -467 -306 -455 -130
rect -421 -306 -409 -130
rect -467 -318 -409 -306
rect -347 -130 -289 -118
rect -347 -306 -335 -130
rect -301 -306 -289 -130
rect -347 -318 -289 -306
rect -89 -130 -31 -118
rect -89 -306 -77 -130
rect -43 -306 -31 -130
rect -89 -318 -31 -306
rect 31 -130 89 -118
rect 31 -306 43 -130
rect 77 -306 89 -130
rect 31 -318 89 -306
rect 289 -130 347 -118
rect 289 -306 301 -130
rect 335 -306 347 -130
rect 289 -318 347 -306
rect 409 -130 467 -118
rect 409 -306 421 -130
rect 455 -306 467 -130
rect 409 -318 467 -306
rect 667 -130 725 -118
rect 667 -306 679 -130
rect 713 -306 725 -130
rect 667 -318 725 -306
rect 787 -130 845 -118
rect 787 -306 799 -130
rect 833 -306 845 -130
rect 787 -318 845 -306
rect 1045 -130 1103 -118
rect 1045 -306 1057 -130
rect 1091 -306 1103 -130
rect 1045 -318 1103 -306
rect 1165 -130 1223 -118
rect 1165 -306 1177 -130
rect 1211 -306 1223 -130
rect 1165 -318 1223 -306
rect 1423 -130 1481 -118
rect 1423 -306 1435 -130
rect 1469 -306 1481 -130
rect 1423 -318 1481 -306
<< mvpdiffc >>
rect -1469 130 -1435 306
rect -1211 130 -1177 306
rect -1091 130 -1057 306
rect -833 130 -799 306
rect -713 130 -679 306
rect -455 130 -421 306
rect -335 130 -301 306
rect -77 130 -43 306
rect 43 130 77 306
rect 301 130 335 306
rect 421 130 455 306
rect 679 130 713 306
rect 799 130 833 306
rect 1057 130 1091 306
rect 1177 130 1211 306
rect 1435 130 1469 306
rect -1469 -306 -1435 -130
rect -1211 -306 -1177 -130
rect -1091 -306 -1057 -130
rect -833 -306 -799 -130
rect -713 -306 -679 -130
rect -455 -306 -421 -130
rect -335 -306 -301 -130
rect -77 -306 -43 -130
rect 43 -306 77 -130
rect 301 -306 335 -130
rect 421 -306 455 -130
rect 679 -306 713 -130
rect 799 -306 833 -130
rect 1057 -306 1091 -130
rect 1177 -306 1211 -130
rect 1435 -306 1469 -130
<< mvnsubdiff >>
rect -1615 537 1615 549
rect -1615 503 -1507 537
rect 1507 503 1615 537
rect -1615 491 1615 503
rect -1615 441 -1557 491
rect -1615 -441 -1603 441
rect -1569 -441 -1557 441
rect 1557 441 1615 491
rect -1615 -491 -1557 -441
rect 1557 -441 1569 441
rect 1603 -441 1615 441
rect 1557 -491 1615 -441
rect -1615 -503 1615 -491
rect -1615 -537 -1507 -503
rect 1507 -537 1615 -503
rect -1615 -549 1615 -537
<< mvnsubdiffcont >>
rect -1507 503 1507 537
rect -1603 -441 -1569 441
rect 1569 -441 1603 441
rect -1507 -537 1507 -503
<< poly >>
rect -1423 399 -1223 415
rect -1423 365 -1407 399
rect -1239 365 -1223 399
rect -1423 318 -1223 365
rect -1045 399 -845 415
rect -1045 365 -1029 399
rect -861 365 -845 399
rect -1045 318 -845 365
rect -667 399 -467 415
rect -667 365 -651 399
rect -483 365 -467 399
rect -667 318 -467 365
rect -289 399 -89 415
rect -289 365 -273 399
rect -105 365 -89 399
rect -289 318 -89 365
rect 89 399 289 415
rect 89 365 105 399
rect 273 365 289 399
rect 89 318 289 365
rect 467 399 667 415
rect 467 365 483 399
rect 651 365 667 399
rect 467 318 667 365
rect 845 399 1045 415
rect 845 365 861 399
rect 1029 365 1045 399
rect 845 318 1045 365
rect 1223 399 1423 415
rect 1223 365 1239 399
rect 1407 365 1423 399
rect 1223 318 1423 365
rect -1423 71 -1223 118
rect -1423 37 -1407 71
rect -1239 37 -1223 71
rect -1423 21 -1223 37
rect -1045 71 -845 118
rect -1045 37 -1029 71
rect -861 37 -845 71
rect -1045 21 -845 37
rect -667 71 -467 118
rect -667 37 -651 71
rect -483 37 -467 71
rect -667 21 -467 37
rect -289 71 -89 118
rect -289 37 -273 71
rect -105 37 -89 71
rect -289 21 -89 37
rect 89 71 289 118
rect 89 37 105 71
rect 273 37 289 71
rect 89 21 289 37
rect 467 71 667 118
rect 467 37 483 71
rect 651 37 667 71
rect 467 21 667 37
rect 845 71 1045 118
rect 845 37 861 71
rect 1029 37 1045 71
rect 845 21 1045 37
rect 1223 71 1423 118
rect 1223 37 1239 71
rect 1407 37 1423 71
rect 1223 21 1423 37
rect -1423 -37 -1223 -21
rect -1423 -71 -1407 -37
rect -1239 -71 -1223 -37
rect -1423 -118 -1223 -71
rect -1045 -37 -845 -21
rect -1045 -71 -1029 -37
rect -861 -71 -845 -37
rect -1045 -118 -845 -71
rect -667 -37 -467 -21
rect -667 -71 -651 -37
rect -483 -71 -467 -37
rect -667 -118 -467 -71
rect -289 -37 -89 -21
rect -289 -71 -273 -37
rect -105 -71 -89 -37
rect -289 -118 -89 -71
rect 89 -37 289 -21
rect 89 -71 105 -37
rect 273 -71 289 -37
rect 89 -118 289 -71
rect 467 -37 667 -21
rect 467 -71 483 -37
rect 651 -71 667 -37
rect 467 -118 667 -71
rect 845 -37 1045 -21
rect 845 -71 861 -37
rect 1029 -71 1045 -37
rect 845 -118 1045 -71
rect 1223 -37 1423 -21
rect 1223 -71 1239 -37
rect 1407 -71 1423 -37
rect 1223 -118 1423 -71
rect -1423 -365 -1223 -318
rect -1423 -399 -1407 -365
rect -1239 -399 -1223 -365
rect -1423 -415 -1223 -399
rect -1045 -365 -845 -318
rect -1045 -399 -1029 -365
rect -861 -399 -845 -365
rect -1045 -415 -845 -399
rect -667 -365 -467 -318
rect -667 -399 -651 -365
rect -483 -399 -467 -365
rect -667 -415 -467 -399
rect -289 -365 -89 -318
rect -289 -399 -273 -365
rect -105 -399 -89 -365
rect -289 -415 -89 -399
rect 89 -365 289 -318
rect 89 -399 105 -365
rect 273 -399 289 -365
rect 89 -415 289 -399
rect 467 -365 667 -318
rect 467 -399 483 -365
rect 651 -399 667 -365
rect 467 -415 667 -399
rect 845 -365 1045 -318
rect 845 -399 861 -365
rect 1029 -399 1045 -365
rect 845 -415 1045 -399
rect 1223 -365 1423 -318
rect 1223 -399 1239 -365
rect 1407 -399 1423 -365
rect 1223 -415 1423 -399
<< polycont >>
rect -1407 365 -1239 399
rect -1029 365 -861 399
rect -651 365 -483 399
rect -273 365 -105 399
rect 105 365 273 399
rect 483 365 651 399
rect 861 365 1029 399
rect 1239 365 1407 399
rect -1407 37 -1239 71
rect -1029 37 -861 71
rect -651 37 -483 71
rect -273 37 -105 71
rect 105 37 273 71
rect 483 37 651 71
rect 861 37 1029 71
rect 1239 37 1407 71
rect -1407 -71 -1239 -37
rect -1029 -71 -861 -37
rect -651 -71 -483 -37
rect -273 -71 -105 -37
rect 105 -71 273 -37
rect 483 -71 651 -37
rect 861 -71 1029 -37
rect 1239 -71 1407 -37
rect -1407 -399 -1239 -365
rect -1029 -399 -861 -365
rect -651 -399 -483 -365
rect -273 -399 -105 -365
rect 105 -399 273 -365
rect 483 -399 651 -365
rect 861 -399 1029 -365
rect 1239 -399 1407 -365
<< locali >>
rect -1603 503 -1507 537
rect 1507 503 1603 537
rect -1603 441 -1569 503
rect 1569 441 1603 503
rect -1423 365 -1407 399
rect -1239 365 -1223 399
rect -1045 365 -1029 399
rect -861 365 -845 399
rect -667 365 -651 399
rect -483 365 -467 399
rect -289 365 -273 399
rect -105 365 -89 399
rect 89 365 105 399
rect 273 365 289 399
rect 467 365 483 399
rect 651 365 667 399
rect 845 365 861 399
rect 1029 365 1045 399
rect 1223 365 1239 399
rect 1407 365 1423 399
rect -1469 306 -1435 322
rect -1469 114 -1435 130
rect -1211 306 -1177 322
rect -1211 114 -1177 130
rect -1091 306 -1057 322
rect -1091 114 -1057 130
rect -833 306 -799 322
rect -833 114 -799 130
rect -713 306 -679 322
rect -713 114 -679 130
rect -455 306 -421 322
rect -455 114 -421 130
rect -335 306 -301 322
rect -335 114 -301 130
rect -77 306 -43 322
rect -77 114 -43 130
rect 43 306 77 322
rect 43 114 77 130
rect 301 306 335 322
rect 301 114 335 130
rect 421 306 455 322
rect 421 114 455 130
rect 679 306 713 322
rect 679 114 713 130
rect 799 306 833 322
rect 799 114 833 130
rect 1057 306 1091 322
rect 1057 114 1091 130
rect 1177 306 1211 322
rect 1177 114 1211 130
rect 1435 306 1469 322
rect 1435 114 1469 130
rect -1423 37 -1407 71
rect -1239 37 -1223 71
rect -1045 37 -1029 71
rect -861 37 -845 71
rect -667 37 -651 71
rect -483 37 -467 71
rect -289 37 -273 71
rect -105 37 -89 71
rect 89 37 105 71
rect 273 37 289 71
rect 467 37 483 71
rect 651 37 667 71
rect 845 37 861 71
rect 1029 37 1045 71
rect 1223 37 1239 71
rect 1407 37 1423 71
rect -1423 -71 -1407 -37
rect -1239 -71 -1223 -37
rect -1045 -71 -1029 -37
rect -861 -71 -845 -37
rect -667 -71 -651 -37
rect -483 -71 -467 -37
rect -289 -71 -273 -37
rect -105 -71 -89 -37
rect 89 -71 105 -37
rect 273 -71 289 -37
rect 467 -71 483 -37
rect 651 -71 667 -37
rect 845 -71 861 -37
rect 1029 -71 1045 -37
rect 1223 -71 1239 -37
rect 1407 -71 1423 -37
rect -1469 -130 -1435 -114
rect -1469 -322 -1435 -306
rect -1211 -130 -1177 -114
rect -1211 -322 -1177 -306
rect -1091 -130 -1057 -114
rect -1091 -322 -1057 -306
rect -833 -130 -799 -114
rect -833 -322 -799 -306
rect -713 -130 -679 -114
rect -713 -322 -679 -306
rect -455 -130 -421 -114
rect -455 -322 -421 -306
rect -335 -130 -301 -114
rect -335 -322 -301 -306
rect -77 -130 -43 -114
rect -77 -322 -43 -306
rect 43 -130 77 -114
rect 43 -322 77 -306
rect 301 -130 335 -114
rect 301 -322 335 -306
rect 421 -130 455 -114
rect 421 -322 455 -306
rect 679 -130 713 -114
rect 679 -322 713 -306
rect 799 -130 833 -114
rect 799 -322 833 -306
rect 1057 -130 1091 -114
rect 1057 -322 1091 -306
rect 1177 -130 1211 -114
rect 1177 -322 1211 -306
rect 1435 -130 1469 -114
rect 1435 -322 1469 -306
rect -1423 -399 -1407 -365
rect -1239 -399 -1223 -365
rect -1045 -399 -1029 -365
rect -861 -399 -845 -365
rect -667 -399 -651 -365
rect -483 -399 -467 -365
rect -289 -399 -273 -365
rect -105 -399 -89 -365
rect 89 -399 105 -365
rect 273 -399 289 -365
rect 467 -399 483 -365
rect 651 -399 667 -365
rect 845 -399 861 -365
rect 1029 -399 1045 -365
rect 1223 -399 1239 -365
rect 1407 -399 1423 -365
rect -1603 -503 -1569 -441
rect 1569 -503 1603 -441
rect -1603 -537 -1507 -503
rect 1507 -537 1603 -503
<< viali >>
rect -1255 503 1255 537
rect -1603 -402 -1569 402
rect -1407 365 -1239 399
rect -1029 365 -861 399
rect -651 365 -483 399
rect -273 365 -105 399
rect 105 365 273 399
rect 483 365 651 399
rect 861 365 1029 399
rect 1239 365 1407 399
rect -1469 130 -1435 306
rect -1211 130 -1177 306
rect -1091 130 -1057 306
rect -833 130 -799 306
rect -713 130 -679 306
rect -455 130 -421 306
rect -335 130 -301 306
rect -77 130 -43 306
rect 43 130 77 306
rect 301 130 335 306
rect 421 130 455 306
rect 679 130 713 306
rect 799 130 833 306
rect 1057 130 1091 306
rect 1177 130 1211 306
rect 1435 130 1469 306
rect -1407 37 -1239 71
rect -1029 37 -861 71
rect -651 37 -483 71
rect -273 37 -105 71
rect 105 37 273 71
rect 483 37 651 71
rect 861 37 1029 71
rect 1239 37 1407 71
rect -1407 -71 -1239 -37
rect -1029 -71 -861 -37
rect -651 -71 -483 -37
rect -273 -71 -105 -37
rect 105 -71 273 -37
rect 483 -71 651 -37
rect 861 -71 1029 -37
rect 1239 -71 1407 -37
rect -1469 -306 -1435 -130
rect -1211 -306 -1177 -130
rect -1091 -306 -1057 -130
rect -833 -306 -799 -130
rect -713 -306 -679 -130
rect -455 -306 -421 -130
rect -335 -306 -301 -130
rect -77 -306 -43 -130
rect 43 -306 77 -130
rect 301 -306 335 -130
rect 421 -306 455 -130
rect 679 -306 713 -130
rect 799 -306 833 -130
rect 1057 -306 1091 -130
rect 1177 -306 1211 -130
rect 1435 -306 1469 -130
rect -1407 -399 -1239 -365
rect -1029 -399 -861 -365
rect -651 -399 -483 -365
rect -273 -399 -105 -365
rect 105 -399 273 -365
rect 483 -399 651 -365
rect 861 -399 1029 -365
rect 1239 -399 1407 -365
rect 1569 -402 1603 402
<< metal1 >>
rect -1267 537 1267 543
rect -1267 503 -1255 537
rect 1255 503 1267 537
rect -1267 497 1267 503
rect -1609 402 -1563 414
rect -1609 -402 -1603 402
rect -1569 -402 -1563 402
rect -1419 399 -1227 405
rect -1419 365 -1407 399
rect -1239 365 -1227 399
rect -1419 359 -1227 365
rect -1041 399 -849 405
rect -1041 365 -1029 399
rect -861 365 -849 399
rect -1041 359 -849 365
rect -663 399 -471 405
rect -663 365 -651 399
rect -483 365 -471 399
rect -663 359 -471 365
rect -285 399 -93 405
rect -285 365 -273 399
rect -105 365 -93 399
rect -285 359 -93 365
rect 93 399 285 405
rect 93 365 105 399
rect 273 365 285 399
rect 93 359 285 365
rect 471 399 663 405
rect 471 365 483 399
rect 651 365 663 399
rect 471 359 663 365
rect 849 399 1041 405
rect 849 365 861 399
rect 1029 365 1041 399
rect 849 359 1041 365
rect 1227 399 1419 405
rect 1227 365 1239 399
rect 1407 365 1419 399
rect 1227 359 1419 365
rect 1563 402 1609 414
rect -1475 306 -1429 318
rect -1475 130 -1469 306
rect -1435 130 -1429 306
rect -1475 118 -1429 130
rect -1217 306 -1171 318
rect -1217 130 -1211 306
rect -1177 130 -1171 306
rect -1217 118 -1171 130
rect -1097 306 -1051 318
rect -1097 130 -1091 306
rect -1057 130 -1051 306
rect -1097 118 -1051 130
rect -839 306 -793 318
rect -839 130 -833 306
rect -799 130 -793 306
rect -839 118 -793 130
rect -719 306 -673 318
rect -719 130 -713 306
rect -679 130 -673 306
rect -719 118 -673 130
rect -461 306 -415 318
rect -461 130 -455 306
rect -421 130 -415 306
rect -461 118 -415 130
rect -341 306 -295 318
rect -341 130 -335 306
rect -301 130 -295 306
rect -341 118 -295 130
rect -83 306 -37 318
rect -83 130 -77 306
rect -43 130 -37 306
rect -83 118 -37 130
rect 37 306 83 318
rect 37 130 43 306
rect 77 130 83 306
rect 37 118 83 130
rect 295 306 341 318
rect 295 130 301 306
rect 335 130 341 306
rect 295 118 341 130
rect 415 306 461 318
rect 415 130 421 306
rect 455 130 461 306
rect 415 118 461 130
rect 673 306 719 318
rect 673 130 679 306
rect 713 130 719 306
rect 673 118 719 130
rect 793 306 839 318
rect 793 130 799 306
rect 833 130 839 306
rect 793 118 839 130
rect 1051 306 1097 318
rect 1051 130 1057 306
rect 1091 130 1097 306
rect 1051 118 1097 130
rect 1171 306 1217 318
rect 1171 130 1177 306
rect 1211 130 1217 306
rect 1171 118 1217 130
rect 1429 306 1475 318
rect 1429 130 1435 306
rect 1469 130 1475 306
rect 1429 118 1475 130
rect -1419 71 -1227 77
rect -1419 37 -1407 71
rect -1239 37 -1227 71
rect -1419 31 -1227 37
rect -1041 71 -849 77
rect -1041 37 -1029 71
rect -861 37 -849 71
rect -1041 31 -849 37
rect -663 71 -471 77
rect -663 37 -651 71
rect -483 37 -471 71
rect -663 31 -471 37
rect -285 71 -93 77
rect -285 37 -273 71
rect -105 37 -93 71
rect -285 31 -93 37
rect 93 71 285 77
rect 93 37 105 71
rect 273 37 285 71
rect 93 31 285 37
rect 471 71 663 77
rect 471 37 483 71
rect 651 37 663 71
rect 471 31 663 37
rect 849 71 1041 77
rect 849 37 861 71
rect 1029 37 1041 71
rect 849 31 1041 37
rect 1227 71 1419 77
rect 1227 37 1239 71
rect 1407 37 1419 71
rect 1227 31 1419 37
rect -1419 -37 -1227 -31
rect -1419 -71 -1407 -37
rect -1239 -71 -1227 -37
rect -1419 -77 -1227 -71
rect -1041 -37 -849 -31
rect -1041 -71 -1029 -37
rect -861 -71 -849 -37
rect -1041 -77 -849 -71
rect -663 -37 -471 -31
rect -663 -71 -651 -37
rect -483 -71 -471 -37
rect -663 -77 -471 -71
rect -285 -37 -93 -31
rect -285 -71 -273 -37
rect -105 -71 -93 -37
rect -285 -77 -93 -71
rect 93 -37 285 -31
rect 93 -71 105 -37
rect 273 -71 285 -37
rect 93 -77 285 -71
rect 471 -37 663 -31
rect 471 -71 483 -37
rect 651 -71 663 -37
rect 471 -77 663 -71
rect 849 -37 1041 -31
rect 849 -71 861 -37
rect 1029 -71 1041 -37
rect 849 -77 1041 -71
rect 1227 -37 1419 -31
rect 1227 -71 1239 -37
rect 1407 -71 1419 -37
rect 1227 -77 1419 -71
rect -1475 -130 -1429 -118
rect -1475 -306 -1469 -130
rect -1435 -306 -1429 -130
rect -1475 -318 -1429 -306
rect -1217 -130 -1171 -118
rect -1217 -306 -1211 -130
rect -1177 -306 -1171 -130
rect -1217 -318 -1171 -306
rect -1097 -130 -1051 -118
rect -1097 -306 -1091 -130
rect -1057 -306 -1051 -130
rect -1097 -318 -1051 -306
rect -839 -130 -793 -118
rect -839 -306 -833 -130
rect -799 -306 -793 -130
rect -839 -318 -793 -306
rect -719 -130 -673 -118
rect -719 -306 -713 -130
rect -679 -306 -673 -130
rect -719 -318 -673 -306
rect -461 -130 -415 -118
rect -461 -306 -455 -130
rect -421 -306 -415 -130
rect -461 -318 -415 -306
rect -341 -130 -295 -118
rect -341 -306 -335 -130
rect -301 -306 -295 -130
rect -341 -318 -295 -306
rect -83 -130 -37 -118
rect -83 -306 -77 -130
rect -43 -306 -37 -130
rect -83 -318 -37 -306
rect 37 -130 83 -118
rect 37 -306 43 -130
rect 77 -306 83 -130
rect 37 -318 83 -306
rect 295 -130 341 -118
rect 295 -306 301 -130
rect 335 -306 341 -130
rect 295 -318 341 -306
rect 415 -130 461 -118
rect 415 -306 421 -130
rect 455 -306 461 -130
rect 415 -318 461 -306
rect 673 -130 719 -118
rect 673 -306 679 -130
rect 713 -306 719 -130
rect 673 -318 719 -306
rect 793 -130 839 -118
rect 793 -306 799 -130
rect 833 -306 839 -130
rect 793 -318 839 -306
rect 1051 -130 1097 -118
rect 1051 -306 1057 -130
rect 1091 -306 1097 -130
rect 1051 -318 1097 -306
rect 1171 -130 1217 -118
rect 1171 -306 1177 -130
rect 1211 -306 1217 -130
rect 1171 -318 1217 -306
rect 1429 -130 1475 -118
rect 1429 -306 1435 -130
rect 1469 -306 1475 -130
rect 1429 -318 1475 -306
rect -1609 -414 -1563 -402
rect -1419 -365 -1227 -359
rect -1419 -399 -1407 -365
rect -1239 -399 -1227 -365
rect -1419 -405 -1227 -399
rect -1041 -365 -849 -359
rect -1041 -399 -1029 -365
rect -861 -399 -849 -365
rect -1041 -405 -849 -399
rect -663 -365 -471 -359
rect -663 -399 -651 -365
rect -483 -399 -471 -365
rect -663 -405 -471 -399
rect -285 -365 -93 -359
rect -285 -399 -273 -365
rect -105 -399 -93 -365
rect -285 -405 -93 -399
rect 93 -365 285 -359
rect 93 -399 105 -365
rect 273 -399 285 -365
rect 93 -405 285 -399
rect 471 -365 663 -359
rect 471 -399 483 -365
rect 651 -399 663 -365
rect 471 -405 663 -399
rect 849 -365 1041 -359
rect 849 -399 861 -365
rect 1029 -399 1041 -365
rect 849 -405 1041 -399
rect 1227 -365 1419 -359
rect 1227 -399 1239 -365
rect 1407 -399 1419 -365
rect 1227 -405 1419 -399
rect 1563 -402 1569 402
rect 1603 -402 1609 402
rect 1563 -414 1609 -402
<< properties >>
string FIXED_BBOX -1586 -520 1586 520
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 2 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 80 viagl 80 viagt 80
string sky130_fd_pr__pfet_g5v0d10v5_U7XX7W parameters
<< end >>
