MACRO tt_um_emilian_rf_playground
  CLASS BLOCK ;
  FOREIGN tt_um_emilian_rf_playground ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.920000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 64.000000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 64.000000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.000000 ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.460400 ;
    ANTENNADIFFAREA 220.414398 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 97.200 205.525 98.010 205.665 ;
        RECT 97.010 205.355 98.010 205.525 ;
      LAYER nwell ;
        RECT 90.205 184.020 91.810 201.860 ;
      LAYER pwell ;
        RECT 92.200 196.465 93.010 201.665 ;
        RECT 93.700 201.525 94.510 201.665 ;
        RECT 93.510 201.355 94.510 201.525 ;
        RECT 92.200 196.295 93.200 196.465 ;
        RECT 92.200 196.155 93.010 196.295 ;
        RECT 93.700 196.155 94.510 201.355 ;
        RECT 92.140 195.475 92.925 195.905 ;
        RECT 93.785 195.425 94.570 195.855 ;
        RECT 93.510 195.260 93.680 195.325 ;
        RECT 92.100 194.425 93.010 195.250 ;
        RECT 93.510 195.155 94.610 195.260 ;
        RECT 92.100 194.320 93.200 194.425 ;
        RECT 93.700 194.330 94.610 195.155 ;
        RECT 93.030 194.255 93.200 194.320 ;
        RECT 93.510 193.910 93.680 193.975 ;
        RECT 92.100 193.075 93.010 193.900 ;
        RECT 93.510 193.805 94.610 193.910 ;
        RECT 92.100 192.970 93.200 193.075 ;
        RECT 93.700 192.980 94.610 193.805 ;
        RECT 93.030 192.905 93.200 192.970 ;
        RECT 93.510 192.560 93.680 192.625 ;
        RECT 92.100 191.725 93.010 192.550 ;
        RECT 93.510 192.455 94.610 192.560 ;
        RECT 92.100 191.620 93.200 191.725 ;
        RECT 93.700 191.630 94.610 192.455 ;
        RECT 93.030 191.555 93.200 191.620 ;
        RECT 93.510 191.210 93.680 191.275 ;
        RECT 92.100 190.375 93.010 191.200 ;
        RECT 93.510 191.105 94.610 191.210 ;
        RECT 92.100 190.270 93.200 190.375 ;
        RECT 93.700 190.280 94.610 191.105 ;
        RECT 93.030 190.205 93.200 190.270 ;
        RECT 93.510 189.860 93.680 189.925 ;
        RECT 92.100 189.025 93.010 189.850 ;
        RECT 93.510 189.755 94.610 189.860 ;
        RECT 92.100 188.920 93.200 189.025 ;
        RECT 93.700 188.930 94.610 189.755 ;
        RECT 93.030 188.855 93.200 188.920 ;
        RECT 93.510 188.510 93.680 188.575 ;
        RECT 92.100 187.675 93.010 188.500 ;
        RECT 93.510 188.405 94.610 188.510 ;
        RECT 92.100 187.570 93.200 187.675 ;
        RECT 93.700 187.580 94.610 188.405 ;
        RECT 93.030 187.505 93.200 187.570 ;
        RECT 93.510 187.160 93.680 187.225 ;
        RECT 92.100 186.325 93.010 187.150 ;
        RECT 93.510 187.055 94.610 187.160 ;
        RECT 92.100 186.220 93.200 186.325 ;
        RECT 93.700 186.230 94.610 187.055 ;
        RECT 93.030 186.155 93.200 186.220 ;
        RECT 93.510 185.810 93.680 185.875 ;
        RECT 92.100 184.975 93.010 185.800 ;
        RECT 93.510 185.705 94.610 185.810 ;
        RECT 92.100 184.870 93.200 184.975 ;
        RECT 93.700 184.880 94.610 185.705 ;
        RECT 93.030 184.805 93.200 184.870 ;
        RECT 92.140 184.225 92.925 184.655 ;
        RECT 93.785 184.225 94.570 184.655 ;
      LAYER nwell ;
        RECT 94.900 184.020 96.505 201.860 ;
      LAYER pwell ;
        RECT 97.200 200.155 98.010 205.355 ;
        RECT 97.010 199.655 97.180 199.825 ;
        RECT 97.200 197.135 97.880 199.560 ;
        RECT 97.285 196.075 98.070 196.505 ;
        RECT 97.200 195.725 97.880 195.865 ;
        RECT 97.010 195.555 97.880 195.725 ;
        RECT 97.200 193.125 97.880 195.555 ;
        RECT 97.200 192.725 97.880 192.865 ;
        RECT 97.010 192.555 97.880 192.725 ;
        RECT 97.200 191.035 97.880 192.555 ;
        RECT 97.200 189.705 97.980 190.765 ;
        RECT 97.010 189.535 97.980 189.705 ;
        RECT 97.200 189.395 97.980 189.535 ;
        RECT 97.285 188.725 98.070 189.155 ;
        RECT 97.200 188.325 98.010 188.465 ;
        RECT 97.010 188.155 98.010 188.325 ;
        RECT 97.200 182.955 98.010 188.155 ;
      LAYER nwell ;
        RECT 98.400 182.760 100.005 205.860 ;
      LAYER pwell ;
        RECT 120.500 200.190 131.400 201.190 ;
        RECT 116.500 199.950 131.400 200.190 ;
        RECT 116.450 196.990 131.400 199.950 ;
        RECT 116.500 196.890 131.400 196.990 ;
      LAYER nwell ;
        RECT 113.810 196.140 120.000 196.150 ;
        RECT 113.800 190.190 120.000 196.140 ;
      LAYER pwell ;
        RECT 120.600 193.490 131.400 196.890 ;
      LAYER nwell ;
        RECT 132.000 194.240 138.200 200.190 ;
        RECT 132.000 194.230 138.190 194.240 ;
      LAYER pwell ;
        RECT 120.600 193.390 135.500 193.490 ;
        RECT 120.600 190.430 135.550 193.390 ;
        RECT 120.600 190.190 135.500 190.430 ;
        RECT 120.600 189.190 131.500 190.190 ;
        RECT 120.500 188.190 131.400 189.190 ;
        RECT 116.500 187.950 131.400 188.190 ;
        RECT 116.450 184.990 131.400 187.950 ;
        RECT 116.500 184.890 131.400 184.990 ;
      LAYER nwell ;
        RECT 113.810 184.140 120.000 184.150 ;
        RECT 113.800 178.190 120.000 184.140 ;
      LAYER pwell ;
        RECT 120.600 181.490 131.400 184.890 ;
      LAYER nwell ;
        RECT 132.000 182.240 138.200 188.190 ;
        RECT 132.000 182.230 138.190 182.240 ;
      LAYER pwell ;
        RECT 120.600 181.390 135.500 181.490 ;
        RECT 120.600 178.430 135.550 181.390 ;
        RECT 120.600 178.190 135.500 178.430 ;
        RECT 120.600 177.190 131.500 178.190 ;
        RECT 120.500 176.190 131.400 177.190 ;
        RECT 116.500 175.950 131.400 176.190 ;
        RECT 116.450 172.990 131.400 175.950 ;
        RECT 116.500 172.890 131.400 172.990 ;
      LAYER nwell ;
        RECT 113.810 172.140 120.000 172.150 ;
        RECT 113.800 166.190 120.000 172.140 ;
      LAYER pwell ;
        RECT 120.600 169.490 131.400 172.890 ;
      LAYER nwell ;
        RECT 132.000 170.240 138.200 176.190 ;
        RECT 132.000 170.230 138.190 170.240 ;
      LAYER pwell ;
        RECT 120.600 169.390 135.500 169.490 ;
        RECT 120.600 166.430 135.550 169.390 ;
        RECT 120.600 166.190 135.500 166.430 ;
        RECT 120.600 165.190 131.500 166.190 ;
        RECT 120.500 164.190 131.400 165.190 ;
        RECT 116.500 163.950 131.400 164.190 ;
        RECT 116.450 160.990 131.400 163.950 ;
        RECT 116.500 160.890 131.400 160.990 ;
      LAYER nwell ;
        RECT 113.810 160.140 120.000 160.150 ;
        RECT 113.800 154.190 120.000 160.140 ;
      LAYER pwell ;
        RECT 120.600 157.490 131.400 160.890 ;
      LAYER nwell ;
        RECT 132.000 158.240 138.200 164.190 ;
        RECT 132.000 158.230 138.190 158.240 ;
      LAYER pwell ;
        RECT 120.600 157.390 135.500 157.490 ;
        RECT 120.600 154.430 135.550 157.390 ;
        RECT 120.600 154.190 135.500 154.430 ;
        RECT 120.600 153.190 131.500 154.190 ;
      LAYER nwell ;
        RECT 123.500 151.200 131.700 151.290 ;
        RECT 120.010 151.090 131.750 151.200 ;
        RECT 120.010 148.290 131.800 151.090 ;
        RECT 120.010 148.240 131.750 148.290 ;
        RECT 112.000 126.000 114.960 132.190 ;
        RECT 108.460 45.250 111.420 51.440 ;
        RECT 113.050 45.180 116.010 51.370 ;
        RECT 118.050 45.000 122.300 63.190 ;
        RECT 124.050 45.000 128.300 63.190 ;
        RECT 130.050 45.000 134.300 63.190 ;
      LAYER pwell ;
        RECT 108.050 33.000 111.010 43.100 ;
        RECT 112.050 33.000 115.010 43.100 ;
        RECT 117.050 33.000 120.010 43.100 ;
        RECT 121.050 33.000 124.010 43.100 ;
        RECT 107.870 13.190 114.700 31.290 ;
        RECT 117.050 13.000 123.880 31.100 ;
        RECT 126.050 25.000 129.010 43.100 ;
        RECT 130.050 25.000 134.300 43.100 ;
        RECT 125.050 22.000 140.870 24.010 ;
        RECT 125.050 19.000 140.870 21.010 ;
        RECT 125.050 14.000 128.010 18.100 ;
        RECT 130.050 14.000 133.010 18.100 ;
      LAYER li1 ;
        RECT 97.010 205.585 97.180 205.670 ;
        RECT 99.730 205.585 99.900 205.670 ;
        RECT 97.010 203.005 98.470 205.585 ;
        RECT 97.010 202.260 97.950 203.005 ;
        RECT 98.640 202.835 99.900 205.585 ;
        RECT 90.310 201.580 90.480 201.670 ;
        RECT 93.030 201.580 93.200 201.670 ;
        RECT 90.310 199.990 90.915 201.580 ;
        RECT 90.310 199.640 92.165 199.990 ;
        RECT 90.310 196.235 90.915 199.640 ;
        RECT 92.485 198.160 93.200 201.580 ;
        RECT 91.655 197.820 93.200 198.160 ;
        RECT 92.485 196.235 93.200 197.820 ;
        RECT 90.310 196.150 90.480 196.235 ;
        RECT 93.030 196.150 93.200 196.235 ;
        RECT 93.510 201.585 93.680 201.670 ;
        RECT 96.230 201.585 96.400 201.670 ;
        RECT 93.510 200.000 94.225 201.585 ;
        RECT 93.510 199.660 95.055 200.000 ;
        RECT 93.510 196.240 94.225 199.660 ;
        RECT 95.795 198.180 96.400 201.585 ;
        RECT 94.545 197.830 96.400 198.180 ;
        RECT 95.795 196.240 96.400 197.830 ;
        RECT 93.510 196.150 93.680 196.240 ;
        RECT 96.230 196.150 96.400 196.240 ;
        RECT 96.855 200.240 97.950 202.260 ;
        RECT 98.120 202.260 99.900 202.835 ;
        RECT 98.120 200.240 100.055 202.260 ;
        RECT 96.855 200.150 97.180 200.240 ;
        RECT 99.730 200.150 100.055 200.240 ;
        RECT 96.855 199.970 97.155 200.150 ;
        RECT 99.755 199.970 100.055 200.150 ;
        RECT 96.855 199.405 97.180 199.970 ;
        RECT 99.730 199.885 100.055 199.970 ;
        RECT 97.820 199.695 98.725 199.865 ;
        RECT 96.855 199.110 97.650 199.405 ;
        RECT 96.855 198.510 97.180 199.110 ;
        RECT 97.820 198.940 97.990 199.695 ;
        RECT 97.375 198.680 97.990 198.940 ;
        RECT 96.855 198.250 97.650 198.510 ;
        RECT 96.855 197.655 97.180 198.250 ;
        RECT 97.820 198.080 97.990 198.680 ;
        RECT 97.375 197.825 97.990 198.080 ;
        RECT 96.855 197.355 97.650 197.655 ;
        RECT 96.855 196.750 97.180 197.355 ;
        RECT 97.820 197.135 97.990 197.825 ;
        RECT 98.160 197.310 98.385 199.525 ;
        RECT 98.555 199.365 98.725 199.695 ;
        RECT 98.895 199.540 100.055 199.885 ;
        RECT 98.555 199.110 99.530 199.365 ;
        RECT 98.555 198.505 98.725 199.110 ;
        RECT 99.730 198.940 100.055 199.540 ;
        RECT 98.895 198.680 100.055 198.940 ;
        RECT 98.555 198.250 99.530 198.505 ;
        RECT 98.555 197.650 98.725 198.250 ;
        RECT 99.730 198.080 100.055 198.680 ;
        RECT 98.895 197.820 100.055 198.080 ;
        RECT 98.555 197.390 99.530 197.650 ;
        RECT 98.555 197.135 98.725 197.390 ;
        RECT 99.730 197.220 100.055 197.820 ;
        RECT 97.820 196.835 98.725 197.135 ;
        RECT 98.895 196.835 100.055 197.220 ;
        RECT 98.155 196.760 98.455 196.835 ;
        RECT 99.730 196.750 100.055 196.835 ;
        RECT 96.855 196.520 97.155 196.750 ;
        RECT 99.755 196.520 100.055 196.750 ;
        RECT 96.855 196.460 97.180 196.520 ;
        RECT 99.730 196.460 100.055 196.520 ;
        RECT 96.855 196.160 97.955 196.460 ;
        RECT 98.555 196.160 100.055 196.460 ;
        RECT 96.855 196.060 97.180 196.160 ;
        RECT 97.360 196.145 97.905 196.160 ;
        RECT 98.565 196.145 99.550 196.160 ;
        RECT 99.730 196.060 100.055 196.160 ;
        RECT 90.310 194.660 90.480 195.920 ;
        RECT 93.030 195.910 93.200 195.920 ;
        RECT 91.155 195.835 91.555 195.860 ;
        RECT 90.660 195.545 91.645 195.835 ;
        RECT 91.155 195.460 91.555 195.545 ;
        RECT 92.305 195.460 94.455 195.910 ;
        RECT 96.855 195.870 97.155 196.060 ;
        RECT 99.755 195.870 100.055 196.060 ;
        RECT 95.355 195.785 95.755 195.860 ;
        RECT 95.065 195.495 96.050 195.785 ;
        RECT 95.355 195.460 95.755 195.495 ;
        RECT 90.650 194.930 92.860 195.160 ;
        RECT 90.650 194.830 91.630 194.930 ;
        RECT 92.230 194.830 92.860 194.930 ;
        RECT 90.310 194.450 91.620 194.660 ;
        RECT 90.310 193.310 90.480 194.450 ;
        RECT 91.800 194.430 92.040 194.760 ;
        RECT 93.030 194.660 93.200 195.460 ;
        RECT 92.210 194.430 93.200 194.660 ;
        RECT 90.650 193.580 92.860 193.810 ;
        RECT 90.650 193.480 91.630 193.580 ;
        RECT 92.230 193.480 92.860 193.580 ;
        RECT 90.310 193.100 91.620 193.310 ;
        RECT 90.310 191.960 90.480 193.100 ;
        RECT 91.800 193.080 92.040 193.410 ;
        RECT 93.030 193.310 93.200 194.430 ;
        RECT 92.210 193.080 93.200 193.310 ;
        RECT 90.650 192.230 92.860 192.460 ;
        RECT 90.650 192.130 91.630 192.230 ;
        RECT 92.230 192.130 92.860 192.230 ;
        RECT 90.310 191.750 91.620 191.960 ;
        RECT 90.310 190.610 90.480 191.750 ;
        RECT 91.800 191.730 92.040 192.060 ;
        RECT 93.030 191.960 93.200 193.080 ;
        RECT 92.210 191.730 93.200 191.960 ;
        RECT 90.650 190.880 92.860 191.110 ;
        RECT 90.650 190.780 91.630 190.880 ;
        RECT 92.230 190.780 92.860 190.880 ;
        RECT 90.310 190.400 91.620 190.610 ;
        RECT 90.310 189.260 90.480 190.400 ;
        RECT 91.800 190.380 92.040 190.710 ;
        RECT 93.030 190.610 93.200 191.730 ;
        RECT 92.210 190.380 93.200 190.610 ;
        RECT 90.650 189.530 92.860 189.760 ;
        RECT 90.650 189.430 91.630 189.530 ;
        RECT 92.230 189.430 92.860 189.530 ;
        RECT 90.310 189.050 91.620 189.260 ;
        RECT 90.310 187.910 90.480 189.050 ;
        RECT 91.800 189.030 92.040 189.360 ;
        RECT 93.030 189.260 93.200 190.380 ;
        RECT 92.210 189.030 93.200 189.260 ;
        RECT 90.650 188.180 92.860 188.410 ;
        RECT 90.650 188.080 91.630 188.180 ;
        RECT 92.230 188.080 92.860 188.180 ;
        RECT 90.310 187.700 91.620 187.910 ;
        RECT 90.310 186.560 90.480 187.700 ;
        RECT 91.800 187.680 92.040 188.010 ;
        RECT 93.030 187.910 93.200 189.030 ;
        RECT 92.210 187.680 93.200 187.910 ;
        RECT 90.650 186.830 92.860 187.060 ;
        RECT 90.650 186.730 91.630 186.830 ;
        RECT 92.230 186.730 92.860 186.830 ;
        RECT 90.310 186.350 91.620 186.560 ;
        RECT 90.310 185.210 90.480 186.350 ;
        RECT 91.800 186.330 92.040 186.660 ;
        RECT 93.030 186.560 93.200 187.680 ;
        RECT 92.210 186.330 93.200 186.560 ;
        RECT 90.650 185.480 92.860 185.710 ;
        RECT 90.650 185.380 91.630 185.480 ;
        RECT 92.230 185.380 92.860 185.480 ;
        RECT 90.310 185.000 91.620 185.210 ;
        RECT 90.310 184.210 90.480 185.000 ;
        RECT 91.800 184.980 92.040 185.310 ;
        RECT 93.030 185.210 93.200 186.330 ;
        RECT 92.210 184.980 93.200 185.210 ;
        RECT 93.030 184.660 93.200 184.980 ;
        RECT 93.510 195.150 93.680 195.460 ;
        RECT 93.510 194.920 94.500 195.150 ;
        RECT 93.510 193.800 93.680 194.920 ;
        RECT 94.670 194.820 94.910 195.150 ;
        RECT 96.230 195.130 96.400 195.870 ;
        RECT 95.090 194.920 96.400 195.130 ;
        RECT 93.850 194.650 94.480 194.750 ;
        RECT 95.080 194.650 96.060 194.750 ;
        RECT 93.850 194.420 96.060 194.650 ;
        RECT 93.510 193.570 94.500 193.800 ;
        RECT 93.510 192.450 93.680 193.570 ;
        RECT 94.670 193.470 94.910 193.800 ;
        RECT 96.230 193.780 96.400 194.920 ;
        RECT 95.090 193.570 96.400 193.780 ;
        RECT 93.850 193.300 94.480 193.400 ;
        RECT 95.080 193.300 96.060 193.400 ;
        RECT 93.850 193.070 96.060 193.300 ;
        RECT 93.510 192.220 94.500 192.450 ;
        RECT 93.510 191.100 93.680 192.220 ;
        RECT 94.670 192.120 94.910 192.450 ;
        RECT 96.230 192.430 96.400 193.570 ;
        RECT 95.090 192.220 96.400 192.430 ;
        RECT 93.850 191.950 94.480 192.050 ;
        RECT 95.080 191.950 96.060 192.050 ;
        RECT 93.850 191.720 96.060 191.950 ;
        RECT 93.510 190.870 94.500 191.100 ;
        RECT 93.510 189.750 93.680 190.870 ;
        RECT 94.670 190.770 94.910 191.100 ;
        RECT 96.230 191.080 96.400 192.220 ;
        RECT 95.090 190.870 96.400 191.080 ;
        RECT 93.850 190.600 94.480 190.700 ;
        RECT 95.080 190.600 96.060 190.700 ;
        RECT 93.850 190.370 96.060 190.600 ;
        RECT 93.510 189.520 94.500 189.750 ;
        RECT 93.510 188.400 93.680 189.520 ;
        RECT 94.670 189.420 94.910 189.750 ;
        RECT 96.230 189.730 96.400 190.870 ;
        RECT 95.090 189.520 96.400 189.730 ;
        RECT 93.850 189.250 94.480 189.350 ;
        RECT 95.080 189.250 96.060 189.350 ;
        RECT 93.850 189.020 96.060 189.250 ;
        RECT 93.510 188.170 94.500 188.400 ;
        RECT 93.510 187.050 93.680 188.170 ;
        RECT 94.670 188.070 94.910 188.400 ;
        RECT 96.230 188.380 96.400 189.520 ;
        RECT 95.090 188.170 96.400 188.380 ;
        RECT 93.850 187.900 94.480 188.000 ;
        RECT 95.080 187.900 96.060 188.000 ;
        RECT 93.850 187.670 96.060 187.900 ;
        RECT 93.510 186.820 94.500 187.050 ;
        RECT 93.510 185.700 93.680 186.820 ;
        RECT 94.670 186.720 94.910 187.050 ;
        RECT 96.230 187.030 96.400 188.170 ;
        RECT 95.090 186.820 96.400 187.030 ;
        RECT 93.850 186.550 94.480 186.650 ;
        RECT 95.080 186.550 96.060 186.650 ;
        RECT 93.850 186.320 96.060 186.550 ;
        RECT 93.510 185.470 94.500 185.700 ;
        RECT 93.510 184.660 93.680 185.470 ;
        RECT 94.670 185.370 94.910 185.700 ;
        RECT 96.230 185.680 96.400 186.820 ;
        RECT 95.090 185.470 96.400 185.680 ;
        RECT 93.850 185.200 94.480 185.300 ;
        RECT 95.080 185.200 96.060 185.300 ;
        RECT 93.850 184.970 96.060 185.200 ;
        RECT 90.660 184.295 91.645 184.585 ;
        RECT 91.155 184.160 91.555 184.295 ;
        RECT 92.305 184.210 94.405 184.660 ;
        RECT 95.065 184.295 96.050 184.585 ;
        RECT 95.455 184.160 95.855 184.295 ;
        RECT 96.230 184.210 96.400 185.470 ;
        RECT 96.855 195.315 97.180 195.870 ;
        RECT 97.350 195.615 99.560 195.785 ;
        RECT 97.350 195.485 97.680 195.615 ;
        RECT 98.590 195.475 99.560 195.615 ;
        RECT 96.855 195.040 97.660 195.315 ;
        RECT 97.850 195.095 98.420 195.445 ;
        RECT 96.855 194.395 97.180 195.040 ;
        RECT 98.590 194.925 98.760 195.475 ;
        RECT 99.730 195.305 100.055 195.870 ;
        RECT 98.930 194.995 100.055 195.305 ;
        RECT 97.440 194.565 98.000 194.860 ;
        RECT 96.855 194.140 97.660 194.395 ;
        RECT 96.855 193.535 97.180 194.140 ;
        RECT 97.830 193.965 98.000 194.565 ;
        RECT 97.440 193.705 98.000 193.965 ;
        RECT 98.170 194.755 98.760 194.925 ;
        RECT 98.170 193.785 98.340 194.755 ;
        RECT 98.930 194.565 99.560 194.825 ;
        RECT 98.930 193.965 99.100 194.565 ;
        RECT 99.730 194.395 100.055 194.995 ;
        RECT 99.270 194.140 100.055 194.395 ;
        RECT 97.830 193.615 98.000 193.705 ;
        RECT 98.510 193.705 99.560 193.965 ;
        RECT 98.510 193.615 98.680 193.705 ;
        RECT 96.855 193.255 97.660 193.535 ;
        RECT 96.855 193.110 97.180 193.255 ;
        RECT 97.830 193.210 98.680 193.615 ;
        RECT 99.730 193.535 100.055 194.140 ;
        RECT 98.860 193.250 100.055 193.535 ;
        RECT 99.730 193.110 100.055 193.250 ;
        RECT 96.855 192.870 97.155 193.110 ;
        RECT 99.755 192.870 100.055 193.110 ;
        RECT 96.855 192.315 97.180 192.870 ;
        RECT 97.350 192.615 99.530 192.785 ;
        RECT 97.350 192.525 97.680 192.615 ;
        RECT 98.590 192.515 99.530 192.615 ;
        RECT 96.855 192.040 97.660 192.315 ;
        RECT 97.840 192.085 98.420 192.445 ;
        RECT 96.855 191.455 97.180 192.040 ;
        RECT 98.590 191.905 98.760 192.515 ;
        RECT 99.730 192.345 100.055 192.870 ;
        RECT 98.950 192.015 100.055 192.345 ;
        RECT 97.350 191.625 97.920 191.830 ;
        RECT 98.090 191.655 98.760 191.905 ;
        RECT 97.750 191.485 97.920 191.625 ;
        RECT 98.950 191.625 99.530 191.810 ;
        RECT 98.950 191.485 99.125 191.625 ;
        RECT 96.855 191.120 97.580 191.455 ;
        RECT 97.750 191.145 99.125 191.485 ;
        RECT 99.730 191.455 100.055 192.015 ;
        RECT 99.305 191.120 100.055 191.455 ;
        RECT 96.855 191.030 97.180 191.120 ;
        RECT 99.730 191.030 100.055 191.120 ;
        RECT 96.855 190.770 97.155 191.030 ;
        RECT 96.855 190.245 97.180 190.770 ;
        RECT 98.155 190.685 98.405 190.810 ;
        RECT 99.755 190.770 100.055 191.030 ;
        RECT 97.350 190.515 99.560 190.685 ;
        RECT 97.350 190.425 97.855 190.515 ;
        RECT 98.655 190.415 99.560 190.515 ;
        RECT 96.855 189.915 97.560 190.245 ;
        RECT 98.155 190.230 98.485 190.345 ;
        RECT 99.730 190.245 100.055 190.770 ;
        RECT 97.730 190.060 98.800 190.230 ;
        RECT 96.855 189.390 97.180 189.915 ;
        RECT 97.730 189.735 97.900 190.060 ;
        RECT 98.155 189.825 98.355 189.860 ;
        RECT 97.350 189.565 97.900 189.735 ;
        RECT 98.080 189.495 98.450 189.825 ;
        RECT 98.630 189.735 98.800 190.060 ;
        RECT 98.970 189.915 100.055 190.245 ;
        RECT 98.630 189.565 99.560 189.735 ;
        RECT 98.155 189.460 98.355 189.495 ;
        RECT 99.730 189.390 100.055 189.915 ;
        RECT 96.855 189.170 97.155 189.390 ;
        RECT 99.755 189.170 100.055 189.390 ;
        RECT 96.855 189.160 97.180 189.170 ;
        RECT 99.730 189.160 100.055 189.170 ;
        RECT 96.855 188.760 97.955 189.160 ;
        RECT 98.555 188.760 100.055 189.160 ;
        RECT 96.855 188.710 97.180 188.760 ;
        RECT 99.730 188.710 100.055 188.760 ;
        RECT 96.855 188.470 97.155 188.710 ;
        RECT 99.755 188.470 100.055 188.710 ;
        RECT 96.855 188.385 97.180 188.470 ;
        RECT 99.730 188.385 100.055 188.470 ;
        RECT 96.855 185.805 98.470 188.385 ;
        RECT 96.855 183.040 97.950 185.805 ;
        RECT 98.640 185.635 100.055 188.385 ;
        RECT 98.120 183.040 100.055 185.635 ;
        RECT 96.855 182.960 97.180 183.040 ;
        RECT 97.010 182.950 97.180 182.960 ;
        RECT 99.730 182.960 100.055 183.040 ;
        RECT 99.730 182.950 99.900 182.960 ;
        RECT 110.100 151.790 112.200 205.790 ;
        RECT 113.000 202.190 139.000 204.190 ;
        RECT 113.000 201.190 114.500 202.190 ;
        RECT 137.500 201.190 139.000 202.190 ;
        RECT 113.000 200.120 114.750 201.190 ;
        RECT 120.500 200.690 131.500 201.190 ;
        RECT 137.250 200.990 139.000 201.190 ;
        RECT 120.500 200.390 127.400 200.690 ;
        RECT 128.100 200.440 129.600 200.690 ;
        RECT 120.500 200.190 121.400 200.390 ;
        RECT 113.000 196.290 116.120 200.120 ;
        RECT 116.500 199.590 121.400 200.190 ;
        RECT 121.930 199.930 123.970 200.100 ;
        RECT 116.500 197.390 116.800 199.590 ;
        RECT 117.480 199.030 119.520 199.200 ;
        RECT 117.140 197.970 117.310 198.970 ;
        RECT 119.690 197.970 119.860 198.970 ;
        RECT 120.100 198.290 121.400 199.590 ;
        RECT 121.590 198.870 121.760 199.870 ;
        RECT 122.400 198.810 123.900 198.890 ;
        RECT 124.140 198.870 124.310 199.870 ;
        RECT 121.930 198.640 123.970 198.810 ;
        RECT 122.400 198.290 123.900 198.640 ;
        RECT 124.600 198.590 127.400 200.390 ;
        RECT 128.030 200.270 130.070 200.440 ;
        RECT 127.690 199.990 127.860 200.210 ;
        RECT 130.240 199.990 130.410 200.210 ;
        RECT 127.690 199.210 130.410 199.990 ;
        RECT 127.700 198.990 130.400 199.210 ;
        RECT 128.030 198.980 130.070 198.990 ;
        RECT 130.600 198.590 131.500 200.690 ;
        RECT 124.600 198.290 131.500 198.590 ;
        RECT 117.480 197.740 119.520 197.910 ;
        RECT 120.100 197.890 131.500 198.290 ;
        RECT 120.100 197.600 127.400 197.890 ;
        RECT 120.100 197.390 121.400 197.600 ;
        RECT 116.500 196.890 121.400 197.390 ;
        RECT 121.950 197.200 123.950 197.340 ;
        RECT 121.930 197.030 123.970 197.200 ;
        RECT 113.000 195.690 119.900 196.290 ;
        RECT 113.000 193.590 114.300 195.690 ;
        RECT 114.885 195.340 118.925 195.400 ;
        RECT 114.600 195.170 119.250 195.340 ;
        RECT 114.500 194.790 119.310 195.170 ;
        RECT 114.500 194.170 114.670 194.790 ;
        RECT 119.140 194.170 119.310 194.790 ;
        RECT 114.885 193.940 118.925 194.110 ;
        RECT 115.100 193.590 118.750 193.940 ;
        RECT 119.600 193.590 119.900 195.690 ;
        RECT 113.000 192.690 119.900 193.590 ;
        RECT 113.000 190.590 114.300 192.690 ;
        RECT 115.100 192.400 118.750 192.690 ;
        RECT 114.885 192.230 118.925 192.400 ;
        RECT 114.500 191.170 114.670 192.170 ;
        RECT 119.140 191.170 119.310 192.170 ;
        RECT 114.885 190.940 118.925 191.110 ;
        RECT 119.600 190.590 119.900 192.690 ;
        RECT 113.000 189.390 119.900 190.590 ;
        RECT 120.500 195.390 121.400 196.890 ;
        RECT 121.590 195.970 121.760 196.970 ;
        RECT 122.400 195.910 123.900 195.990 ;
        RECT 124.140 195.970 124.310 196.970 ;
        RECT 121.930 195.740 123.970 195.910 ;
        RECT 122.400 195.390 123.900 195.740 ;
        RECT 124.600 195.690 127.400 197.600 ;
        RECT 128.100 197.540 129.600 197.890 ;
        RECT 128.030 197.370 130.070 197.540 ;
        RECT 127.690 197.090 127.860 197.310 ;
        RECT 130.240 197.090 130.410 197.310 ;
        RECT 127.690 196.310 130.410 197.090 ;
        RECT 127.700 196.090 130.400 196.310 ;
        RECT 128.030 196.080 130.070 196.090 ;
        RECT 130.600 195.690 131.500 197.890 ;
        RECT 124.600 195.390 131.500 195.690 ;
        RECT 120.500 194.990 131.500 195.390 ;
        RECT 120.500 194.690 127.400 194.990 ;
        RECT 120.500 192.490 121.400 194.690 ;
        RECT 121.930 194.290 123.970 194.300 ;
        RECT 121.600 194.070 124.300 194.290 ;
        RECT 121.590 193.290 124.310 194.070 ;
        RECT 121.590 193.070 121.760 193.290 ;
        RECT 124.140 193.070 124.310 193.290 ;
        RECT 121.930 192.840 123.970 193.010 ;
        RECT 122.400 192.490 123.900 192.840 ;
        RECT 124.600 192.780 127.400 194.690 ;
        RECT 128.100 194.640 129.600 194.990 ;
        RECT 128.030 194.470 130.070 194.640 ;
        RECT 127.690 193.410 127.860 194.410 ;
        RECT 128.100 194.390 129.600 194.470 ;
        RECT 130.240 193.410 130.410 194.410 ;
        RECT 130.600 193.490 131.500 194.990 ;
        RECT 132.100 199.790 139.000 200.990 ;
        RECT 132.100 197.690 132.400 199.790 ;
        RECT 133.075 199.270 137.115 199.440 ;
        RECT 132.690 198.210 132.860 199.210 ;
        RECT 137.330 198.210 137.500 199.210 ;
        RECT 133.075 197.980 137.115 198.150 ;
        RECT 133.250 197.690 136.900 197.980 ;
        RECT 137.700 197.690 139.000 199.790 ;
        RECT 132.100 196.790 139.000 197.690 ;
        RECT 132.100 194.690 132.400 196.790 ;
        RECT 133.250 196.440 136.900 196.790 ;
        RECT 133.075 196.270 137.115 196.440 ;
        RECT 132.690 195.590 132.860 196.210 ;
        RECT 137.330 195.590 137.500 196.210 ;
        RECT 132.690 195.210 137.500 195.590 ;
        RECT 132.750 195.040 137.400 195.210 ;
        RECT 133.075 194.980 137.115 195.040 ;
        RECT 137.700 194.690 139.000 196.790 ;
        RECT 132.100 194.090 139.000 194.690 ;
        RECT 128.030 193.180 130.070 193.350 ;
        RECT 128.050 193.040 130.050 193.180 ;
        RECT 130.600 192.990 135.500 193.490 ;
        RECT 130.600 192.780 131.900 192.990 ;
        RECT 124.600 192.490 131.900 192.780 ;
        RECT 120.500 192.090 131.900 192.490 ;
        RECT 132.480 192.470 134.520 192.640 ;
        RECT 120.500 191.790 127.400 192.090 ;
        RECT 120.500 189.690 121.400 191.790 ;
        RECT 121.930 191.390 123.970 191.400 ;
        RECT 121.600 191.170 124.300 191.390 ;
        RECT 121.590 190.390 124.310 191.170 ;
        RECT 121.590 190.170 121.760 190.390 ;
        RECT 124.140 190.170 124.310 190.390 ;
        RECT 121.930 189.940 123.970 190.110 ;
        RECT 124.600 189.990 127.400 191.790 ;
        RECT 128.100 191.740 129.600 192.090 ;
        RECT 128.030 191.570 130.070 191.740 ;
        RECT 127.690 190.510 127.860 191.510 ;
        RECT 128.100 191.490 129.600 191.570 ;
        RECT 130.240 190.510 130.410 191.510 ;
        RECT 130.600 190.790 131.900 192.090 ;
        RECT 132.140 191.410 132.310 192.410 ;
        RECT 134.690 191.410 134.860 192.410 ;
        RECT 132.480 191.180 134.520 191.350 ;
        RECT 135.200 190.790 135.500 192.990 ;
        RECT 128.030 190.280 130.070 190.450 ;
        RECT 130.600 190.190 135.500 190.790 ;
        RECT 135.880 190.260 139.000 194.090 ;
        RECT 130.600 189.990 131.500 190.190 ;
        RECT 122.400 189.690 123.900 189.940 ;
        RECT 124.600 189.690 131.500 189.990 ;
        RECT 113.000 188.120 114.750 189.390 ;
        RECT 120.500 188.690 131.500 189.690 ;
        RECT 137.250 188.990 139.000 190.260 ;
        RECT 120.500 188.390 127.400 188.690 ;
        RECT 128.100 188.440 129.600 188.690 ;
        RECT 120.500 188.190 121.400 188.390 ;
        RECT 113.000 184.290 116.120 188.120 ;
        RECT 116.500 187.590 121.400 188.190 ;
        RECT 121.930 187.930 123.970 188.100 ;
        RECT 116.500 185.390 116.800 187.590 ;
        RECT 117.480 187.030 119.520 187.200 ;
        RECT 117.140 185.970 117.310 186.970 ;
        RECT 119.690 185.970 119.860 186.970 ;
        RECT 120.100 186.290 121.400 187.590 ;
        RECT 121.590 186.870 121.760 187.870 ;
        RECT 122.400 186.810 123.900 186.890 ;
        RECT 124.140 186.870 124.310 187.870 ;
        RECT 121.930 186.640 123.970 186.810 ;
        RECT 122.400 186.290 123.900 186.640 ;
        RECT 124.600 186.590 127.400 188.390 ;
        RECT 128.030 188.270 130.070 188.440 ;
        RECT 127.690 187.990 127.860 188.210 ;
        RECT 130.240 187.990 130.410 188.210 ;
        RECT 127.690 187.210 130.410 187.990 ;
        RECT 127.700 186.990 130.400 187.210 ;
        RECT 128.030 186.980 130.070 186.990 ;
        RECT 130.600 186.590 131.500 188.690 ;
        RECT 124.600 186.290 131.500 186.590 ;
        RECT 117.480 185.740 119.520 185.910 ;
        RECT 120.100 185.890 131.500 186.290 ;
        RECT 120.100 185.600 127.400 185.890 ;
        RECT 120.100 185.390 121.400 185.600 ;
        RECT 116.500 184.890 121.400 185.390 ;
        RECT 121.950 185.200 123.950 185.340 ;
        RECT 121.930 185.030 123.970 185.200 ;
        RECT 113.000 183.690 119.900 184.290 ;
        RECT 113.000 181.590 114.300 183.690 ;
        RECT 114.885 183.340 118.925 183.400 ;
        RECT 114.600 183.170 119.250 183.340 ;
        RECT 114.500 182.790 119.310 183.170 ;
        RECT 114.500 182.170 114.670 182.790 ;
        RECT 119.140 182.170 119.310 182.790 ;
        RECT 114.885 181.940 118.925 182.110 ;
        RECT 115.100 181.590 118.750 181.940 ;
        RECT 119.600 181.590 119.900 183.690 ;
        RECT 113.000 180.690 119.900 181.590 ;
        RECT 113.000 178.590 114.300 180.690 ;
        RECT 115.100 180.400 118.750 180.690 ;
        RECT 114.885 180.230 118.925 180.400 ;
        RECT 114.500 179.170 114.670 180.170 ;
        RECT 119.140 179.170 119.310 180.170 ;
        RECT 114.885 178.940 118.925 179.110 ;
        RECT 119.600 178.590 119.900 180.690 ;
        RECT 113.000 177.390 119.900 178.590 ;
        RECT 120.500 183.390 121.400 184.890 ;
        RECT 121.590 183.970 121.760 184.970 ;
        RECT 122.400 183.910 123.900 183.990 ;
        RECT 124.140 183.970 124.310 184.970 ;
        RECT 121.930 183.740 123.970 183.910 ;
        RECT 122.400 183.390 123.900 183.740 ;
        RECT 124.600 183.690 127.400 185.600 ;
        RECT 128.100 185.540 129.600 185.890 ;
        RECT 128.030 185.370 130.070 185.540 ;
        RECT 127.690 185.090 127.860 185.310 ;
        RECT 130.240 185.090 130.410 185.310 ;
        RECT 127.690 184.310 130.410 185.090 ;
        RECT 127.700 184.090 130.400 184.310 ;
        RECT 128.030 184.080 130.070 184.090 ;
        RECT 130.600 183.690 131.500 185.890 ;
        RECT 124.600 183.390 131.500 183.690 ;
        RECT 120.500 182.990 131.500 183.390 ;
        RECT 120.500 182.690 127.400 182.990 ;
        RECT 120.500 180.490 121.400 182.690 ;
        RECT 121.930 182.290 123.970 182.300 ;
        RECT 121.600 182.070 124.300 182.290 ;
        RECT 121.590 181.290 124.310 182.070 ;
        RECT 121.590 181.070 121.760 181.290 ;
        RECT 124.140 181.070 124.310 181.290 ;
        RECT 121.930 180.840 123.970 181.010 ;
        RECT 122.400 180.490 123.900 180.840 ;
        RECT 124.600 180.780 127.400 182.690 ;
        RECT 128.100 182.640 129.600 182.990 ;
        RECT 128.030 182.470 130.070 182.640 ;
        RECT 127.690 181.410 127.860 182.410 ;
        RECT 128.100 182.390 129.600 182.470 ;
        RECT 130.240 181.410 130.410 182.410 ;
        RECT 130.600 181.490 131.500 182.990 ;
        RECT 132.100 187.790 139.000 188.990 ;
        RECT 132.100 185.690 132.400 187.790 ;
        RECT 133.075 187.270 137.115 187.440 ;
        RECT 132.690 186.210 132.860 187.210 ;
        RECT 137.330 186.210 137.500 187.210 ;
        RECT 133.075 185.980 137.115 186.150 ;
        RECT 133.250 185.690 136.900 185.980 ;
        RECT 137.700 185.690 139.000 187.790 ;
        RECT 132.100 184.790 139.000 185.690 ;
        RECT 132.100 182.690 132.400 184.790 ;
        RECT 133.250 184.440 136.900 184.790 ;
        RECT 133.075 184.270 137.115 184.440 ;
        RECT 132.690 183.590 132.860 184.210 ;
        RECT 137.330 183.590 137.500 184.210 ;
        RECT 132.690 183.210 137.500 183.590 ;
        RECT 132.750 183.040 137.400 183.210 ;
        RECT 133.075 182.980 137.115 183.040 ;
        RECT 137.700 182.690 139.000 184.790 ;
        RECT 132.100 182.090 139.000 182.690 ;
        RECT 128.030 181.180 130.070 181.350 ;
        RECT 128.050 181.040 130.050 181.180 ;
        RECT 130.600 180.990 135.500 181.490 ;
        RECT 130.600 180.780 131.900 180.990 ;
        RECT 124.600 180.490 131.900 180.780 ;
        RECT 120.500 180.090 131.900 180.490 ;
        RECT 132.480 180.470 134.520 180.640 ;
        RECT 120.500 179.790 127.400 180.090 ;
        RECT 120.500 177.690 121.400 179.790 ;
        RECT 121.930 179.390 123.970 179.400 ;
        RECT 121.600 179.170 124.300 179.390 ;
        RECT 121.590 178.390 124.310 179.170 ;
        RECT 121.590 178.170 121.760 178.390 ;
        RECT 124.140 178.170 124.310 178.390 ;
        RECT 121.930 177.940 123.970 178.110 ;
        RECT 124.600 177.990 127.400 179.790 ;
        RECT 128.100 179.740 129.600 180.090 ;
        RECT 128.030 179.570 130.070 179.740 ;
        RECT 127.690 178.510 127.860 179.510 ;
        RECT 128.100 179.490 129.600 179.570 ;
        RECT 130.240 178.510 130.410 179.510 ;
        RECT 130.600 178.790 131.900 180.090 ;
        RECT 132.140 179.410 132.310 180.410 ;
        RECT 134.690 179.410 134.860 180.410 ;
        RECT 132.480 179.180 134.520 179.350 ;
        RECT 135.200 178.790 135.500 180.990 ;
        RECT 128.030 178.280 130.070 178.450 ;
        RECT 130.600 178.190 135.500 178.790 ;
        RECT 135.880 178.260 139.000 182.090 ;
        RECT 130.600 177.990 131.500 178.190 ;
        RECT 122.400 177.690 123.900 177.940 ;
        RECT 124.600 177.690 131.500 177.990 ;
        RECT 113.000 176.120 114.750 177.390 ;
        RECT 120.500 176.690 131.500 177.690 ;
        RECT 137.250 176.990 139.000 178.260 ;
        RECT 120.500 176.390 127.400 176.690 ;
        RECT 128.100 176.440 129.600 176.690 ;
        RECT 120.500 176.190 121.400 176.390 ;
        RECT 113.000 172.290 116.120 176.120 ;
        RECT 116.500 175.590 121.400 176.190 ;
        RECT 121.930 175.930 123.970 176.100 ;
        RECT 116.500 173.390 116.800 175.590 ;
        RECT 117.480 175.030 119.520 175.200 ;
        RECT 117.140 173.970 117.310 174.970 ;
        RECT 119.690 173.970 119.860 174.970 ;
        RECT 120.100 174.290 121.400 175.590 ;
        RECT 121.590 174.870 121.760 175.870 ;
        RECT 122.400 174.810 123.900 174.890 ;
        RECT 124.140 174.870 124.310 175.870 ;
        RECT 121.930 174.640 123.970 174.810 ;
        RECT 122.400 174.290 123.900 174.640 ;
        RECT 124.600 174.590 127.400 176.390 ;
        RECT 128.030 176.270 130.070 176.440 ;
        RECT 127.690 175.990 127.860 176.210 ;
        RECT 130.240 175.990 130.410 176.210 ;
        RECT 127.690 175.210 130.410 175.990 ;
        RECT 127.700 174.990 130.400 175.210 ;
        RECT 128.030 174.980 130.070 174.990 ;
        RECT 130.600 174.590 131.500 176.690 ;
        RECT 124.600 174.290 131.500 174.590 ;
        RECT 117.480 173.740 119.520 173.910 ;
        RECT 120.100 173.890 131.500 174.290 ;
        RECT 120.100 173.600 127.400 173.890 ;
        RECT 120.100 173.390 121.400 173.600 ;
        RECT 116.500 172.890 121.400 173.390 ;
        RECT 121.950 173.200 123.950 173.340 ;
        RECT 121.930 173.030 123.970 173.200 ;
        RECT 113.000 171.690 119.900 172.290 ;
        RECT 113.000 169.590 114.300 171.690 ;
        RECT 114.885 171.340 118.925 171.400 ;
        RECT 114.600 171.170 119.250 171.340 ;
        RECT 114.500 170.790 119.310 171.170 ;
        RECT 114.500 170.170 114.670 170.790 ;
        RECT 119.140 170.170 119.310 170.790 ;
        RECT 114.885 169.940 118.925 170.110 ;
        RECT 115.100 169.590 118.750 169.940 ;
        RECT 119.600 169.590 119.900 171.690 ;
        RECT 113.000 168.690 119.900 169.590 ;
        RECT 113.000 166.590 114.300 168.690 ;
        RECT 115.100 168.400 118.750 168.690 ;
        RECT 114.885 168.230 118.925 168.400 ;
        RECT 114.500 167.170 114.670 168.170 ;
        RECT 119.140 167.170 119.310 168.170 ;
        RECT 114.885 166.940 118.925 167.110 ;
        RECT 119.600 166.590 119.900 168.690 ;
        RECT 113.000 165.390 119.900 166.590 ;
        RECT 120.500 171.390 121.400 172.890 ;
        RECT 121.590 171.970 121.760 172.970 ;
        RECT 122.400 171.910 123.900 171.990 ;
        RECT 124.140 171.970 124.310 172.970 ;
        RECT 121.930 171.740 123.970 171.910 ;
        RECT 122.400 171.390 123.900 171.740 ;
        RECT 124.600 171.690 127.400 173.600 ;
        RECT 128.100 173.540 129.600 173.890 ;
        RECT 128.030 173.370 130.070 173.540 ;
        RECT 127.690 173.090 127.860 173.310 ;
        RECT 130.240 173.090 130.410 173.310 ;
        RECT 127.690 172.310 130.410 173.090 ;
        RECT 127.700 172.090 130.400 172.310 ;
        RECT 128.030 172.080 130.070 172.090 ;
        RECT 130.600 171.690 131.500 173.890 ;
        RECT 124.600 171.390 131.500 171.690 ;
        RECT 120.500 170.990 131.500 171.390 ;
        RECT 120.500 170.690 127.400 170.990 ;
        RECT 120.500 168.490 121.400 170.690 ;
        RECT 121.930 170.290 123.970 170.300 ;
        RECT 121.600 170.070 124.300 170.290 ;
        RECT 121.590 169.290 124.310 170.070 ;
        RECT 121.590 169.070 121.760 169.290 ;
        RECT 124.140 169.070 124.310 169.290 ;
        RECT 121.930 168.840 123.970 169.010 ;
        RECT 122.400 168.490 123.900 168.840 ;
        RECT 124.600 168.780 127.400 170.690 ;
        RECT 128.100 170.640 129.600 170.990 ;
        RECT 128.030 170.470 130.070 170.640 ;
        RECT 127.690 169.410 127.860 170.410 ;
        RECT 128.100 170.390 129.600 170.470 ;
        RECT 130.240 169.410 130.410 170.410 ;
        RECT 130.600 169.490 131.500 170.990 ;
        RECT 132.100 175.790 139.000 176.990 ;
        RECT 132.100 173.690 132.400 175.790 ;
        RECT 133.075 175.270 137.115 175.440 ;
        RECT 132.690 174.210 132.860 175.210 ;
        RECT 137.330 174.210 137.500 175.210 ;
        RECT 133.075 173.980 137.115 174.150 ;
        RECT 133.250 173.690 136.900 173.980 ;
        RECT 137.700 173.690 139.000 175.790 ;
        RECT 132.100 172.790 139.000 173.690 ;
        RECT 132.100 170.690 132.400 172.790 ;
        RECT 133.250 172.440 136.900 172.790 ;
        RECT 133.075 172.270 137.115 172.440 ;
        RECT 132.690 171.590 132.860 172.210 ;
        RECT 137.330 171.590 137.500 172.210 ;
        RECT 132.690 171.210 137.500 171.590 ;
        RECT 132.750 171.040 137.400 171.210 ;
        RECT 133.075 170.980 137.115 171.040 ;
        RECT 137.700 170.690 139.000 172.790 ;
        RECT 132.100 170.090 139.000 170.690 ;
        RECT 128.030 169.180 130.070 169.350 ;
        RECT 128.050 169.040 130.050 169.180 ;
        RECT 130.600 168.990 135.500 169.490 ;
        RECT 130.600 168.780 131.900 168.990 ;
        RECT 124.600 168.490 131.900 168.780 ;
        RECT 120.500 168.090 131.900 168.490 ;
        RECT 132.480 168.470 134.520 168.640 ;
        RECT 120.500 167.790 127.400 168.090 ;
        RECT 120.500 165.690 121.400 167.790 ;
        RECT 121.930 167.390 123.970 167.400 ;
        RECT 121.600 167.170 124.300 167.390 ;
        RECT 121.590 166.390 124.310 167.170 ;
        RECT 121.590 166.170 121.760 166.390 ;
        RECT 124.140 166.170 124.310 166.390 ;
        RECT 121.930 165.940 123.970 166.110 ;
        RECT 124.600 165.990 127.400 167.790 ;
        RECT 128.100 167.740 129.600 168.090 ;
        RECT 128.030 167.570 130.070 167.740 ;
        RECT 127.690 166.510 127.860 167.510 ;
        RECT 128.100 167.490 129.600 167.570 ;
        RECT 130.240 166.510 130.410 167.510 ;
        RECT 130.600 166.790 131.900 168.090 ;
        RECT 132.140 167.410 132.310 168.410 ;
        RECT 134.690 167.410 134.860 168.410 ;
        RECT 132.480 167.180 134.520 167.350 ;
        RECT 135.200 166.790 135.500 168.990 ;
        RECT 128.030 166.280 130.070 166.450 ;
        RECT 130.600 166.190 135.500 166.790 ;
        RECT 135.880 166.260 139.000 170.090 ;
        RECT 130.600 165.990 131.500 166.190 ;
        RECT 122.400 165.690 123.900 165.940 ;
        RECT 124.600 165.690 131.500 165.990 ;
        RECT 113.000 164.120 114.750 165.390 ;
        RECT 120.500 164.690 131.500 165.690 ;
        RECT 137.250 164.990 139.000 166.260 ;
        RECT 120.500 164.390 127.400 164.690 ;
        RECT 128.100 164.440 129.600 164.690 ;
        RECT 120.500 164.190 121.400 164.390 ;
        RECT 113.000 160.290 116.120 164.120 ;
        RECT 116.500 163.590 121.400 164.190 ;
        RECT 121.930 163.930 123.970 164.100 ;
        RECT 116.500 161.390 116.800 163.590 ;
        RECT 117.480 163.030 119.520 163.200 ;
        RECT 117.140 161.970 117.310 162.970 ;
        RECT 119.690 161.970 119.860 162.970 ;
        RECT 120.100 162.290 121.400 163.590 ;
        RECT 121.590 162.870 121.760 163.870 ;
        RECT 122.400 162.810 123.900 162.890 ;
        RECT 124.140 162.870 124.310 163.870 ;
        RECT 121.930 162.640 123.970 162.810 ;
        RECT 122.400 162.290 123.900 162.640 ;
        RECT 124.600 162.590 127.400 164.390 ;
        RECT 128.030 164.270 130.070 164.440 ;
        RECT 127.690 163.990 127.860 164.210 ;
        RECT 130.240 163.990 130.410 164.210 ;
        RECT 127.690 163.210 130.410 163.990 ;
        RECT 127.700 162.990 130.400 163.210 ;
        RECT 128.030 162.980 130.070 162.990 ;
        RECT 130.600 162.590 131.500 164.690 ;
        RECT 124.600 162.290 131.500 162.590 ;
        RECT 117.480 161.740 119.520 161.910 ;
        RECT 120.100 161.890 131.500 162.290 ;
        RECT 120.100 161.600 127.400 161.890 ;
        RECT 120.100 161.390 121.400 161.600 ;
        RECT 116.500 160.890 121.400 161.390 ;
        RECT 121.950 161.200 123.950 161.340 ;
        RECT 121.930 161.030 123.970 161.200 ;
        RECT 113.000 159.690 119.900 160.290 ;
        RECT 113.000 157.590 114.300 159.690 ;
        RECT 114.885 159.340 118.925 159.400 ;
        RECT 114.600 159.170 119.250 159.340 ;
        RECT 114.500 158.790 119.310 159.170 ;
        RECT 114.500 158.170 114.670 158.790 ;
        RECT 119.140 158.170 119.310 158.790 ;
        RECT 114.885 157.940 118.925 158.110 ;
        RECT 115.100 157.590 118.750 157.940 ;
        RECT 119.600 157.590 119.900 159.690 ;
        RECT 113.000 156.690 119.900 157.590 ;
        RECT 113.000 154.590 114.300 156.690 ;
        RECT 115.100 156.400 118.750 156.690 ;
        RECT 114.885 156.230 118.925 156.400 ;
        RECT 114.500 155.170 114.670 156.170 ;
        RECT 119.140 155.170 119.310 156.170 ;
        RECT 114.885 154.940 118.925 155.110 ;
        RECT 119.600 154.590 119.900 156.690 ;
        RECT 113.000 153.690 119.900 154.590 ;
        RECT 120.500 159.390 121.400 160.890 ;
        RECT 121.590 159.970 121.760 160.970 ;
        RECT 122.400 159.910 123.900 159.990 ;
        RECT 124.140 159.970 124.310 160.970 ;
        RECT 121.930 159.740 123.970 159.910 ;
        RECT 122.400 159.390 123.900 159.740 ;
        RECT 124.600 159.690 127.400 161.600 ;
        RECT 128.100 161.540 129.600 161.890 ;
        RECT 128.030 161.370 130.070 161.540 ;
        RECT 127.690 161.090 127.860 161.310 ;
        RECT 130.240 161.090 130.410 161.310 ;
        RECT 127.690 160.310 130.410 161.090 ;
        RECT 127.700 160.090 130.400 160.310 ;
        RECT 128.030 160.080 130.070 160.090 ;
        RECT 130.600 159.690 131.500 161.890 ;
        RECT 124.600 159.390 131.500 159.690 ;
        RECT 120.500 158.990 131.500 159.390 ;
        RECT 120.500 158.690 127.400 158.990 ;
        RECT 120.500 156.490 121.400 158.690 ;
        RECT 121.930 158.290 123.970 158.300 ;
        RECT 121.600 158.070 124.300 158.290 ;
        RECT 121.590 157.290 124.310 158.070 ;
        RECT 121.590 157.070 121.760 157.290 ;
        RECT 124.140 157.070 124.310 157.290 ;
        RECT 121.930 156.840 123.970 157.010 ;
        RECT 122.400 156.490 123.900 156.840 ;
        RECT 124.600 156.780 127.400 158.690 ;
        RECT 128.100 158.640 129.600 158.990 ;
        RECT 128.030 158.470 130.070 158.640 ;
        RECT 127.690 157.410 127.860 158.410 ;
        RECT 128.100 158.390 129.600 158.470 ;
        RECT 130.240 157.410 130.410 158.410 ;
        RECT 130.600 157.490 131.500 158.990 ;
        RECT 132.100 163.790 139.000 164.990 ;
        RECT 132.100 161.690 132.400 163.790 ;
        RECT 133.075 163.270 137.115 163.440 ;
        RECT 132.690 162.210 132.860 163.210 ;
        RECT 137.330 162.210 137.500 163.210 ;
        RECT 133.075 161.980 137.115 162.150 ;
        RECT 133.250 161.690 136.900 161.980 ;
        RECT 137.700 161.690 139.000 163.790 ;
        RECT 132.100 160.790 139.000 161.690 ;
        RECT 132.100 158.690 132.400 160.790 ;
        RECT 133.250 160.440 136.900 160.790 ;
        RECT 133.075 160.270 137.115 160.440 ;
        RECT 132.690 159.590 132.860 160.210 ;
        RECT 137.330 159.590 137.500 160.210 ;
        RECT 132.690 159.210 137.500 159.590 ;
        RECT 132.750 159.040 137.400 159.210 ;
        RECT 133.075 158.980 137.115 159.040 ;
        RECT 137.700 158.690 139.000 160.790 ;
        RECT 132.100 158.090 139.000 158.690 ;
        RECT 128.030 157.180 130.070 157.350 ;
        RECT 128.050 157.040 130.050 157.180 ;
        RECT 130.600 156.990 135.500 157.490 ;
        RECT 130.600 156.780 131.900 156.990 ;
        RECT 124.600 156.490 131.900 156.780 ;
        RECT 120.500 156.090 131.900 156.490 ;
        RECT 132.480 156.470 134.520 156.640 ;
        RECT 120.500 155.790 127.400 156.090 ;
        RECT 120.500 153.690 121.400 155.790 ;
        RECT 121.930 155.390 123.970 155.400 ;
        RECT 121.600 155.170 124.300 155.390 ;
        RECT 121.590 154.390 124.310 155.170 ;
        RECT 121.590 154.170 121.760 154.390 ;
        RECT 124.140 154.170 124.310 154.390 ;
        RECT 121.930 153.940 123.970 154.110 ;
        RECT 124.600 153.990 127.400 155.790 ;
        RECT 128.100 155.740 129.600 156.090 ;
        RECT 128.030 155.570 130.070 155.740 ;
        RECT 127.690 154.510 127.860 155.510 ;
        RECT 128.100 155.490 129.600 155.570 ;
        RECT 130.240 154.510 130.410 155.510 ;
        RECT 130.600 154.790 131.900 156.090 ;
        RECT 132.140 155.410 132.310 156.410 ;
        RECT 134.690 155.410 134.860 156.410 ;
        RECT 132.480 155.180 134.520 155.350 ;
        RECT 135.200 154.790 135.500 156.990 ;
        RECT 128.030 154.280 130.070 154.450 ;
        RECT 130.600 154.190 135.500 154.790 ;
        RECT 135.880 154.260 139.000 158.090 ;
        RECT 130.600 153.990 131.500 154.190 ;
        RECT 122.400 153.690 123.900 153.940 ;
        RECT 124.600 153.690 131.500 153.990 ;
        RECT 113.000 152.190 120.000 153.690 ;
        RECT 120.500 152.690 131.500 153.690 ;
        RECT 137.250 153.190 139.000 154.260 ;
        RECT 137.255 152.690 139.000 153.190 ;
        RECT 139.500 152.690 142.500 203.890 ;
        RECT 113.000 152.090 119.900 152.190 ;
        RECT 112.900 151.790 119.900 152.090 ;
        RECT 110.100 151.290 119.900 151.790 ;
        RECT 120.500 151.690 135.300 152.690 ;
        RECT 110.100 151.090 131.700 151.290 ;
        RECT 110.100 150.850 131.800 151.090 ;
        RECT 110.100 149.690 120.400 150.850 ;
        RECT 123.500 150.790 131.800 150.850 ;
        RECT 121.100 150.450 125.000 150.490 ;
        RECT 121.085 150.280 125.125 150.450 ;
        RECT 110.000 148.690 120.400 149.690 ;
        RECT 120.700 149.220 120.870 150.220 ;
        RECT 121.100 149.790 125.000 150.280 ;
        RECT 125.340 149.220 125.510 150.220 ;
        RECT 121.600 149.160 124.700 149.190 ;
        RECT 121.085 148.990 125.125 149.160 ;
        RECT 121.600 148.690 124.700 148.990 ;
        RECT 125.740 148.690 126.020 150.790 ;
        RECT 126.635 150.280 130.675 150.450 ;
        RECT 126.250 149.220 126.420 150.220 ;
        RECT 130.890 149.220 131.060 150.220 ;
        RECT 126.800 149.160 130.500 149.190 ;
        RECT 126.635 148.990 130.675 149.160 ;
        RECT 126.800 148.690 130.500 148.990 ;
        RECT 131.300 148.690 131.800 150.790 ;
        RECT 132.400 149.490 135.300 151.690 ;
        RECT 137.255 151.190 142.500 152.690 ;
        RECT 137.500 148.690 142.500 151.190 ;
        RECT 110.000 146.890 142.500 148.690 ;
        RECT 110.000 146.190 126.400 146.890 ;
        RECT 130.300 146.190 142.500 146.890 ;
        RECT 112.000 132.010 112.800 132.100 ;
        RECT 112.000 131.840 114.780 132.010 ;
        RECT 112.000 131.115 112.800 131.840 ;
        RECT 112.980 131.330 114.200 131.500 ;
        RECT 113.100 131.115 114.200 131.330 ;
        RECT 112.000 127.075 112.920 131.115 ;
        RECT 113.100 127.075 114.210 131.115 ;
        RECT 112.000 126.350 112.800 127.075 ;
        RECT 113.100 126.860 114.200 127.075 ;
        RECT 112.980 126.690 114.200 126.860 ;
        RECT 113.100 126.650 114.200 126.690 ;
        RECT 114.610 126.350 114.780 131.840 ;
        RECT 112.000 126.200 114.780 126.350 ;
        RECT 112.180 126.180 114.780 126.200 ;
        RECT 105.050 62.840 143.050 67.000 ;
        RECT 105.050 62.115 118.850 62.840 ;
        RECT 119.030 62.330 120.030 62.500 ;
        RECT 120.320 62.330 121.320 62.500 ;
        RECT 121.500 62.115 124.800 62.840 ;
        RECT 125.030 62.330 126.030 62.500 ;
        RECT 126.320 62.330 127.320 62.500 ;
        RECT 127.550 62.115 130.800 62.840 ;
        RECT 131.030 62.330 132.030 62.500 ;
        RECT 132.320 62.330 133.320 62.500 ;
        RECT 133.550 62.115 143.050 62.840 ;
        RECT 105.050 51.090 118.970 62.115 ;
        RECT 105.050 45.600 108.810 51.090 ;
        RECT 111.070 51.000 118.970 51.090 ;
        RECT 109.150 50.750 109.750 50.800 ;
        RECT 109.150 50.580 110.440 50.750 ;
        RECT 111.070 50.700 113.950 51.000 ;
        RECT 111.070 50.680 114.350 50.700 ;
        RECT 109.150 46.110 109.750 50.580 ;
        RECT 111.070 50.510 115.030 50.680 ;
        RECT 110.500 49.850 110.670 50.365 ;
        RECT 111.070 49.850 114.350 50.510 ;
        RECT 110.500 46.700 114.350 49.850 ;
        RECT 110.500 46.325 110.670 46.700 ;
        RECT 109.150 45.940 110.440 46.110 ;
        RECT 109.150 45.900 109.750 45.940 ;
        RECT 111.070 45.600 113.050 46.700 ;
        RECT 105.050 45.400 113.050 45.600 ;
        RECT 113.230 45.530 113.400 46.700 ;
        RECT 113.750 46.040 114.350 46.700 ;
        RECT 115.090 46.255 115.260 50.295 ;
        RECT 113.750 45.870 115.030 46.040 ;
        RECT 113.750 45.800 114.350 45.870 ;
        RECT 115.660 45.530 115.830 51.000 ;
        RECT 113.230 45.400 115.830 45.530 ;
        RECT 116.050 46.075 118.970 51.000 ;
        RECT 120.090 46.075 120.260 62.115 ;
        RECT 121.380 61.850 124.970 62.115 ;
        RECT 121.350 46.450 124.970 61.850 ;
        RECT 121.380 46.075 124.970 46.450 ;
        RECT 126.090 46.075 126.260 62.115 ;
        RECT 127.380 46.075 130.970 62.115 ;
        RECT 132.090 46.075 132.260 62.115 ;
        RECT 133.380 46.400 143.050 62.115 ;
        RECT 133.380 46.075 137.000 46.400 ;
        RECT 116.050 45.400 118.850 46.075 ;
        RECT 119.030 45.690 120.030 45.860 ;
        RECT 120.320 45.690 121.320 45.860 ;
        RECT 105.050 45.350 118.850 45.400 ;
        RECT 121.500 45.350 124.800 46.075 ;
        RECT 125.030 45.690 126.030 45.860 ;
        RECT 126.320 45.690 127.320 45.860 ;
        RECT 127.550 45.350 130.800 46.075 ;
        RECT 131.030 45.690 132.030 45.860 ;
        RECT 132.320 45.690 133.320 45.860 ;
        RECT 133.550 45.350 137.000 46.075 ;
        RECT 105.050 45.000 137.000 45.350 ;
        RECT 105.050 42.700 137.050 43.200 ;
        RECT 105.050 42.500 108.650 42.700 ;
        RECT 110.450 42.500 112.400 42.700 ;
        RECT 105.050 33.350 108.400 42.500 ;
        RECT 109.030 42.240 110.030 42.410 ;
        RECT 108.800 34.030 108.970 42.070 ;
        RECT 110.090 34.030 110.260 42.070 ;
        RECT 109.030 33.690 110.030 33.860 ;
        RECT 110.660 33.350 112.400 42.500 ;
        RECT 113.030 42.240 114.030 42.410 ;
        RECT 112.800 34.030 112.970 42.070 ;
        RECT 114.090 34.030 114.260 42.070 ;
        RECT 113.030 33.690 114.030 33.860 ;
        RECT 114.650 33.350 117.400 42.700 ;
        RECT 118.030 42.240 119.030 42.410 ;
        RECT 117.800 34.030 117.970 42.070 ;
        RECT 119.090 34.030 119.260 42.070 ;
        RECT 118.030 33.690 119.030 33.860 ;
        RECT 119.660 33.350 121.400 42.700 ;
        RECT 122.030 42.240 123.030 42.410 ;
        RECT 121.800 34.030 121.970 42.070 ;
        RECT 123.090 34.030 123.260 42.070 ;
        RECT 122.030 33.690 123.030 33.860 ;
        RECT 123.650 33.350 126.400 42.700 ;
        RECT 127.030 42.400 128.030 42.410 ;
        RECT 105.050 30.900 126.400 33.350 ;
        RECT 105.050 13.550 108.250 30.900 ;
        RECT 114.250 30.650 126.400 30.900 ;
        RECT 108.850 30.430 109.850 30.600 ;
        RECT 110.140 30.430 111.140 30.600 ;
        RECT 111.430 30.430 112.430 30.600 ;
        RECT 112.720 30.430 113.720 30.600 ;
        RECT 108.620 14.220 108.790 30.260 ;
        RECT 109.910 14.220 110.080 30.260 ;
        RECT 111.200 14.220 111.370 30.260 ;
        RECT 112.490 14.220 112.660 30.260 ;
        RECT 113.780 14.220 113.950 30.260 ;
        RECT 108.850 13.880 109.850 14.050 ;
        RECT 110.140 13.880 111.140 14.050 ;
        RECT 111.430 13.880 112.430 14.050 ;
        RECT 112.720 13.880 113.720 14.050 ;
        RECT 114.250 13.550 117.550 30.650 ;
        RECT 118.030 30.240 119.030 30.410 ;
        RECT 119.320 30.240 120.320 30.410 ;
        RECT 120.610 30.240 121.610 30.410 ;
        RECT 121.900 30.240 122.900 30.410 ;
        RECT 117.800 14.030 117.970 30.070 ;
        RECT 119.090 14.030 119.260 30.070 ;
        RECT 120.380 14.030 120.550 30.070 ;
        RECT 121.670 14.030 121.840 30.070 ;
        RECT 122.960 14.030 123.130 30.070 ;
        RECT 123.530 25.350 126.400 30.650 ;
        RECT 126.650 42.240 128.030 42.400 ;
        RECT 126.650 25.860 127.650 42.240 ;
        RECT 128.250 42.070 130.850 42.700 ;
        RECT 131.030 42.240 132.030 42.410 ;
        RECT 132.320 42.240 133.320 42.410 ;
        RECT 133.550 42.070 137.000 42.700 ;
        RECT 128.090 26.030 130.970 42.070 ;
        RECT 132.090 26.030 132.260 42.070 ;
        RECT 133.380 26.050 137.000 42.070 ;
        RECT 133.380 26.030 138.600 26.050 ;
        RECT 126.650 25.690 128.030 25.860 ;
        RECT 126.650 25.600 127.650 25.690 ;
        RECT 128.250 25.350 130.850 26.030 ;
        RECT 133.550 25.950 138.600 26.030 ;
        RECT 131.030 25.690 132.030 25.860 ;
        RECT 132.320 25.690 133.320 25.860 ;
        RECT 133.550 25.350 143.050 25.950 ;
        RECT 123.530 23.600 143.050 25.350 ;
        RECT 123.530 22.400 125.400 23.600 ;
        RECT 125.880 22.830 128.040 23.180 ;
        RECT 137.880 22.830 140.040 23.180 ;
        RECT 140.450 22.400 143.050 23.600 ;
        RECT 123.530 20.650 143.050 22.400 ;
        RECT 123.530 19.350 125.400 20.650 ;
        RECT 125.880 19.830 128.040 20.180 ;
        RECT 137.880 19.830 140.040 20.180 ;
        RECT 140.450 19.350 143.050 20.650 ;
        RECT 123.530 17.750 143.050 19.350 ;
        RECT 123.530 14.400 125.450 17.750 ;
        RECT 127.550 17.700 143.050 17.750 ;
        RECT 126.030 17.240 127.030 17.410 ;
        RECT 125.800 15.030 125.970 17.070 ;
        RECT 127.090 16.950 127.260 17.070 ;
        RECT 127.550 16.950 130.450 17.700 ;
        RECT 131.100 17.410 131.950 17.500 ;
        RECT 132.350 17.450 143.050 17.700 ;
        RECT 131.030 17.240 132.030 17.410 ;
        RECT 131.100 17.200 131.950 17.240 ;
        RECT 131.200 17.150 131.900 17.200 ;
        RECT 127.090 15.110 130.450 16.950 ;
        RECT 127.090 15.030 127.260 15.110 ;
        RECT 126.030 14.690 127.030 14.860 ;
        RECT 127.550 14.400 130.450 15.110 ;
        RECT 130.800 16.450 130.970 17.070 ;
        RECT 131.550 16.450 131.900 17.150 ;
        RECT 130.800 15.450 131.900 16.450 ;
        RECT 130.800 15.030 130.970 15.450 ;
        RECT 131.550 14.950 131.900 15.450 ;
        RECT 132.090 16.900 132.260 17.070 ;
        RECT 132.660 16.900 143.050 17.450 ;
        RECT 132.090 15.200 143.050 16.900 ;
        RECT 132.090 15.030 132.260 15.200 ;
        RECT 131.200 14.900 131.900 14.950 ;
        RECT 131.100 14.860 131.950 14.900 ;
        RECT 131.030 14.690 132.030 14.860 ;
        RECT 132.660 14.700 143.050 15.200 ;
        RECT 131.100 14.600 131.950 14.690 ;
        RECT 132.500 14.550 143.050 14.700 ;
        RECT 123.530 14.350 130.700 14.400 ;
        RECT 132.350 14.350 143.050 14.550 ;
        RECT 118.030 13.690 119.030 13.860 ;
        RECT 119.320 13.690 120.320 13.860 ;
        RECT 120.610 13.690 121.610 13.860 ;
        RECT 121.900 13.690 122.900 13.860 ;
        RECT 105.050 13.350 117.550 13.550 ;
        RECT 123.530 13.350 143.050 14.350 ;
        RECT 105.050 10.000 143.050 13.350 ;
      LAYER met1 ;
        RECT 98.600 207.650 99.500 208.300 ;
        RECT 83.000 205.550 83.700 205.580 ;
        RECT 90.155 205.550 90.855 205.760 ;
        RECT 96.055 205.670 97.055 205.690 ;
        RECT 96.055 205.660 97.335 205.670 ;
        RECT 83.000 204.850 90.855 205.550 ;
        RECT 83.000 204.820 83.700 204.850 ;
        RECT 90.155 197.710 90.855 204.850 ;
        RECT 92.875 201.660 93.835 201.670 ;
        RECT 91.175 201.310 91.535 201.610 ;
        RECT 90.155 196.210 90.955 197.710 ;
        RECT 90.155 184.060 90.655 196.210 ;
        RECT 91.205 195.920 91.505 201.310 ;
        RECT 91.125 195.860 91.585 195.920 ;
        RECT 90.855 195.460 91.585 195.860 ;
        RECT 90.955 195.400 91.585 195.460 ;
        RECT 90.955 184.620 91.255 195.400 ;
        RECT 91.755 195.190 92.155 195.410 ;
        RECT 91.480 194.900 92.350 195.190 ;
        RECT 91.840 194.710 92.070 194.740 ;
        RECT 91.805 193.840 92.105 194.710 ;
        RECT 91.480 193.550 92.350 193.840 ;
        RECT 91.840 193.360 92.070 193.390 ;
        RECT 91.805 192.490 92.105 193.360 ;
        RECT 91.480 192.200 92.350 192.490 ;
        RECT 91.840 191.960 92.070 192.040 ;
        RECT 91.805 191.140 92.105 191.960 ;
        RECT 91.480 190.850 92.350 191.140 ;
        RECT 91.840 190.660 92.070 190.690 ;
        RECT 91.805 189.790 92.105 190.660 ;
        RECT 91.480 189.500 92.350 189.790 ;
        RECT 91.840 189.310 92.070 189.340 ;
        RECT 91.805 188.440 92.105 189.310 ;
        RECT 91.480 188.150 92.350 188.440 ;
        RECT 91.840 187.960 92.070 187.990 ;
        RECT 91.805 187.090 92.105 187.960 ;
        RECT 91.480 186.800 92.350 187.090 ;
        RECT 91.840 186.610 92.070 186.640 ;
        RECT 91.805 185.740 92.105 186.610 ;
        RECT 91.480 185.450 92.350 185.740 ;
        RECT 91.755 184.760 92.155 185.310 ;
        RECT 90.955 184.560 91.585 184.620 ;
        RECT 90.855 184.160 91.585 184.560 ;
        RECT 91.125 184.100 91.585 184.160 ;
        RECT 92.855 184.060 93.855 201.660 ;
        RECT 94.455 201.360 95.155 205.660 ;
        RECT 96.055 204.630 97.355 205.660 ;
        RECT 96.075 201.660 96.555 201.670 ;
        RECT 95.505 201.610 95.805 201.640 ;
        RECT 95.455 201.280 95.805 201.610 ;
        RECT 95.455 195.920 95.755 201.280 ;
        RECT 96.055 197.710 96.555 201.660 ;
        RECT 95.955 196.210 96.555 197.710 ;
        RECT 95.325 195.860 95.785 195.920 ;
        RECT 95.155 195.460 95.855 195.860 ;
        RECT 94.555 194.860 94.955 195.460 ;
        RECT 95.325 195.400 95.785 195.460 ;
        RECT 94.640 194.840 94.870 194.860 ;
        RECT 94.360 194.390 95.230 194.680 ;
        RECT 94.605 193.510 94.905 194.390 ;
        RECT 94.640 193.490 94.870 193.510 ;
        RECT 94.360 193.040 95.230 193.330 ;
        RECT 94.605 192.160 94.905 193.040 ;
        RECT 94.640 192.140 94.870 192.160 ;
        RECT 94.360 191.690 95.230 191.980 ;
        RECT 94.605 190.810 94.905 191.690 ;
        RECT 94.640 190.790 94.870 190.810 ;
        RECT 94.360 190.340 95.230 190.630 ;
        RECT 94.555 189.810 94.905 190.340 ;
        RECT 94.605 189.460 94.905 189.810 ;
        RECT 94.640 189.440 94.870 189.460 ;
        RECT 94.360 188.990 95.230 189.280 ;
        RECT 94.605 188.110 94.905 188.990 ;
        RECT 94.640 188.090 94.870 188.110 ;
        RECT 94.360 187.640 95.230 187.930 ;
        RECT 94.605 186.760 94.905 187.640 ;
        RECT 94.640 186.740 94.870 186.760 ;
        RECT 94.360 186.290 95.230 186.580 ;
        RECT 94.605 185.410 94.905 186.290 ;
        RECT 94.640 185.390 94.870 185.410 ;
        RECT 94.360 184.940 95.230 185.230 ;
        RECT 94.605 184.710 95.005 184.940 ;
        RECT 95.455 184.620 95.755 195.400 ;
        RECT 95.425 184.560 95.885 184.620 ;
        RECT 95.155 184.160 95.885 184.560 ;
        RECT 95.425 184.100 95.885 184.160 ;
        RECT 96.055 184.060 96.555 196.210 ;
        RECT 96.855 182.960 97.355 204.630 ;
        RECT 98.055 197.760 98.455 206.930 ;
        RECT 97.655 197.560 98.455 197.760 ;
        RECT 97.655 197.510 98.405 197.560 ;
        RECT 97.655 193.460 97.905 197.510 ;
        RECT 98.855 197.160 99.255 207.650 ;
        RECT 99.575 205.660 100.055 205.670 ;
        RECT 98.155 197.120 99.255 197.160 ;
        RECT 98.125 196.760 99.255 197.120 ;
        RECT 98.125 196.700 98.485 196.760 ;
        RECT 98.075 195.410 98.385 195.470 ;
        RECT 98.075 195.160 99.155 195.410 ;
        RECT 98.075 195.100 98.385 195.160 ;
        RECT 98.075 193.460 98.385 193.520 ;
        RECT 97.655 193.210 98.405 193.460 ;
        RECT 98.075 193.150 98.385 193.210 ;
        RECT 98.125 192.050 98.435 192.420 ;
        RECT 98.155 190.870 98.405 192.050 ;
        RECT 98.905 191.470 99.155 195.160 ;
        RECT 98.825 191.110 99.155 191.470 ;
        RECT 98.825 191.100 99.135 191.110 ;
        RECT 98.125 190.500 98.435 190.870 ;
        RECT 98.125 189.860 98.385 189.920 ;
        RECT 98.055 189.360 98.555 189.860 ;
        RECT 99.555 182.960 100.055 205.660 ;
        RECT 96.855 182.950 97.335 182.960 ;
        RECT 99.575 182.950 100.055 182.960 ;
        RECT 110.100 151.790 112.200 205.790 ;
        RECT 113.000 202.190 139.000 204.190 ;
        RECT 113.000 201.190 114.500 202.190 ;
        RECT 137.500 201.190 139.000 202.190 ;
        RECT 113.000 200.120 114.750 201.190 ;
        RECT 120.500 200.690 131.400 201.190 ;
        RECT 137.250 200.990 139.000 201.190 ;
        RECT 120.500 200.440 127.400 200.690 ;
        RECT 128.100 200.470 129.600 200.690 ;
        RECT 120.500 200.390 121.450 200.440 ;
        RECT 120.500 200.190 121.400 200.390 ;
        RECT 113.000 196.290 116.120 200.120 ;
        RECT 116.500 199.590 121.400 200.190 ;
        RECT 122.000 200.130 123.950 200.240 ;
        RECT 121.950 199.900 123.950 200.130 ;
        RECT 116.500 197.390 116.800 199.590 ;
        RECT 117.700 199.230 119.500 199.390 ;
        RECT 117.500 199.000 119.500 199.230 ;
        RECT 117.110 198.840 117.340 198.950 ;
        RECT 117.700 198.940 119.500 199.000 ;
        RECT 117.700 198.840 119.250 198.940 ;
        RECT 117.100 198.790 117.400 198.840 ;
        RECT 119.660 198.790 119.890 198.950 ;
        RECT 117.100 198.690 117.500 198.790 ;
        RECT 119.500 198.690 119.900 198.790 ;
        RECT 117.100 198.240 119.900 198.690 ;
        RECT 117.100 198.090 117.500 198.240 ;
        RECT 119.550 198.090 119.900 198.240 ;
        RECT 120.100 198.290 121.400 199.590 ;
        RECT 121.560 199.690 121.790 199.850 ;
        RECT 124.110 199.690 124.340 199.850 ;
        RECT 121.560 199.090 124.340 199.690 ;
        RECT 121.560 198.890 121.790 199.090 ;
        RECT 124.110 198.890 124.340 199.090 ;
        RECT 122.400 198.840 123.900 198.890 ;
        RECT 121.950 198.610 123.950 198.840 ;
        RECT 122.400 198.290 123.900 198.610 ;
        RECT 124.600 198.590 127.400 200.440 ;
        RECT 128.050 200.240 130.050 200.470 ;
        RECT 127.660 199.990 127.890 200.190 ;
        RECT 130.210 200.180 130.440 200.190 ;
        RECT 130.210 200.040 130.500 200.180 ;
        RECT 130.100 199.990 130.500 200.040 ;
        RECT 127.660 199.230 130.500 199.990 ;
        RECT 127.700 199.040 130.500 199.230 ;
        RECT 127.700 198.990 130.400 199.040 ;
        RECT 128.050 198.950 130.050 198.990 ;
        RECT 130.700 198.590 131.400 200.690 ;
        RECT 124.600 198.290 131.400 198.590 ;
        RECT 117.100 198.040 117.400 198.090 ;
        RECT 117.110 197.990 117.340 198.040 ;
        RECT 119.660 197.990 119.890 198.090 ;
        RECT 117.800 197.940 119.400 197.990 ;
        RECT 117.500 197.710 119.500 197.940 ;
        RECT 120.100 197.890 131.400 198.290 ;
        RECT 117.800 197.540 119.450 197.710 ;
        RECT 120.100 197.690 127.400 197.890 ;
        RECT 120.100 197.390 121.400 197.690 ;
        RECT 124.550 197.640 127.400 197.690 ;
        RECT 122.000 197.490 122.500 197.540 ;
        RECT 116.500 196.890 121.400 197.390 ;
        RECT 121.950 197.000 123.950 197.490 ;
        RECT 113.000 195.720 119.900 196.290 ;
        RECT 113.000 193.990 114.300 195.720 ;
        RECT 119.580 195.690 119.900 195.720 ;
        RECT 114.905 195.390 118.905 195.430 ;
        RECT 114.500 195.150 119.300 195.390 ;
        RECT 114.470 194.290 119.340 195.150 ;
        RECT 114.470 194.190 114.700 194.290 ;
        RECT 119.110 194.190 119.340 194.290 ;
        RECT 114.905 193.990 118.905 194.140 ;
        RECT 119.600 193.990 119.900 195.690 ;
        RECT 113.000 192.390 119.900 193.990 ;
        RECT 113.000 192.290 118.905 192.390 ;
        RECT 113.000 190.590 114.300 192.290 ;
        RECT 114.905 192.200 118.905 192.290 ;
        RECT 114.470 191.990 114.700 192.150 ;
        RECT 119.110 191.990 119.340 192.150 ;
        RECT 114.470 191.490 119.340 191.990 ;
        RECT 114.470 191.390 114.800 191.490 ;
        RECT 114.470 191.190 114.700 191.390 ;
        RECT 115.600 191.340 115.900 191.490 ;
        RECT 119.100 191.390 119.340 191.490 ;
        RECT 116.900 191.140 118.700 191.240 ;
        RECT 119.110 191.190 119.340 191.390 ;
        RECT 114.905 190.910 118.905 191.140 ;
        RECT 116.900 190.740 118.700 190.910 ;
        RECT 119.600 190.590 119.900 192.390 ;
        RECT 113.000 189.390 119.900 190.590 ;
        RECT 120.600 195.390 121.400 196.890 ;
        RECT 121.560 196.790 121.790 196.950 ;
        RECT 124.110 196.790 124.340 196.950 ;
        RECT 121.560 196.190 124.340 196.790 ;
        RECT 121.560 195.990 121.790 196.190 ;
        RECT 124.110 195.990 124.340 196.190 ;
        RECT 122.400 195.940 123.900 195.990 ;
        RECT 121.950 195.710 123.950 195.940 ;
        RECT 122.400 195.390 123.900 195.710 ;
        RECT 124.600 195.690 127.400 197.640 ;
        RECT 128.100 197.570 129.600 197.890 ;
        RECT 128.050 197.340 130.050 197.570 ;
        RECT 127.660 197.090 127.890 197.290 ;
        RECT 130.210 197.090 130.440 197.290 ;
        RECT 127.660 196.330 130.440 197.090 ;
        RECT 127.700 196.090 130.400 196.330 ;
        RECT 128.050 196.050 130.050 196.090 ;
        RECT 130.600 195.690 131.400 197.890 ;
        RECT 124.600 195.390 131.400 195.690 ;
        RECT 120.600 194.990 131.400 195.390 ;
        RECT 120.600 194.690 127.400 194.990 ;
        RECT 120.600 192.490 121.400 194.690 ;
        RECT 121.950 194.290 123.950 194.330 ;
        RECT 121.600 194.050 124.300 194.290 ;
        RECT 121.560 193.290 124.340 194.050 ;
        RECT 121.560 193.090 121.790 193.290 ;
        RECT 124.110 193.090 124.340 193.290 ;
        RECT 121.950 192.810 123.950 193.040 ;
        RECT 122.400 192.490 123.900 192.810 ;
        RECT 124.600 192.740 127.400 194.690 ;
        RECT 128.100 194.670 129.600 194.990 ;
        RECT 128.050 194.440 130.050 194.670 ;
        RECT 128.100 194.390 129.600 194.440 ;
        RECT 127.660 194.190 127.890 194.390 ;
        RECT 130.210 194.190 130.440 194.390 ;
        RECT 127.660 193.590 130.440 194.190 ;
        RECT 127.660 193.430 127.890 193.590 ;
        RECT 130.210 193.430 130.440 193.590 ;
        RECT 130.600 193.490 131.400 194.990 ;
        RECT 132.100 199.790 139.000 200.990 ;
        RECT 132.100 197.990 132.400 199.790 ;
        RECT 133.300 199.470 135.100 199.640 ;
        RECT 133.095 199.240 137.095 199.470 ;
        RECT 132.660 198.990 132.890 199.190 ;
        RECT 133.300 199.140 135.100 199.240 ;
        RECT 132.660 198.890 132.900 198.990 ;
        RECT 136.100 198.890 136.400 199.040 ;
        RECT 137.300 198.990 137.530 199.190 ;
        RECT 137.200 198.890 137.530 198.990 ;
        RECT 132.660 198.390 137.530 198.890 ;
        RECT 132.660 198.230 132.890 198.390 ;
        RECT 137.300 198.230 137.530 198.390 ;
        RECT 133.095 198.090 137.095 198.180 ;
        RECT 137.700 198.090 139.000 199.790 ;
        RECT 133.095 197.990 139.000 198.090 ;
        RECT 132.100 196.390 139.000 197.990 ;
        RECT 132.100 194.690 132.400 196.390 ;
        RECT 133.095 196.240 137.095 196.390 ;
        RECT 132.660 196.090 132.890 196.190 ;
        RECT 137.300 196.090 137.530 196.190 ;
        RECT 132.660 195.230 137.530 196.090 ;
        RECT 132.700 194.990 137.500 195.230 ;
        RECT 133.095 194.950 137.095 194.990 ;
        RECT 132.100 194.660 132.420 194.690 ;
        RECT 137.700 194.660 139.000 196.390 ;
        RECT 132.100 194.090 139.000 194.660 ;
        RECT 128.050 192.890 130.050 193.380 ;
        RECT 130.600 192.990 135.500 193.490 ;
        RECT 129.500 192.840 130.000 192.890 ;
        RECT 124.600 192.690 127.450 192.740 ;
        RECT 130.600 192.690 131.900 192.990 ;
        RECT 124.600 192.490 131.900 192.690 ;
        RECT 132.550 192.670 134.200 192.840 ;
        RECT 120.600 192.090 131.900 192.490 ;
        RECT 132.500 192.440 134.500 192.670 ;
        RECT 132.600 192.390 134.200 192.440 ;
        RECT 132.110 192.290 132.340 192.390 ;
        RECT 134.660 192.340 134.890 192.390 ;
        RECT 134.600 192.290 134.900 192.340 ;
        RECT 120.600 191.790 127.400 192.090 ;
        RECT 120.600 189.690 121.300 191.790 ;
        RECT 121.950 191.390 123.950 191.430 ;
        RECT 121.600 191.340 124.300 191.390 ;
        RECT 121.500 191.150 124.300 191.340 ;
        RECT 121.500 190.390 124.340 191.150 ;
        RECT 121.500 190.340 121.900 190.390 ;
        RECT 121.500 190.200 121.790 190.340 ;
        RECT 121.560 190.190 121.790 190.200 ;
        RECT 124.110 190.190 124.340 190.390 ;
        RECT 121.950 189.910 123.950 190.140 ;
        RECT 124.600 189.940 127.400 191.790 ;
        RECT 128.100 191.770 129.600 192.090 ;
        RECT 128.050 191.540 130.050 191.770 ;
        RECT 128.100 191.490 129.600 191.540 ;
        RECT 127.660 191.290 127.890 191.490 ;
        RECT 130.210 191.290 130.440 191.490 ;
        RECT 127.660 190.690 130.440 191.290 ;
        RECT 127.660 190.530 127.890 190.690 ;
        RECT 130.210 190.530 130.440 190.690 ;
        RECT 130.600 190.790 131.900 192.090 ;
        RECT 132.100 192.140 132.450 192.290 ;
        RECT 134.500 192.140 134.900 192.290 ;
        RECT 132.100 191.690 134.900 192.140 ;
        RECT 132.100 191.590 132.500 191.690 ;
        RECT 134.500 191.590 134.900 191.690 ;
        RECT 132.110 191.430 132.340 191.590 ;
        RECT 134.600 191.540 134.900 191.590 ;
        RECT 132.750 191.440 134.300 191.540 ;
        RECT 132.500 191.380 134.300 191.440 ;
        RECT 134.660 191.430 134.890 191.540 ;
        RECT 132.500 191.150 134.500 191.380 ;
        RECT 132.500 190.990 134.300 191.150 ;
        RECT 135.200 190.790 135.500 192.990 ;
        RECT 128.050 190.250 130.050 190.480 ;
        RECT 128.050 190.140 130.000 190.250 ;
        RECT 130.600 190.190 135.500 190.790 ;
        RECT 135.880 190.260 139.000 194.090 ;
        RECT 130.600 189.990 131.500 190.190 ;
        RECT 130.550 189.940 131.500 189.990 ;
        RECT 122.400 189.690 123.900 189.910 ;
        RECT 124.600 189.690 131.500 189.940 ;
        RECT 113.000 188.120 114.750 189.390 ;
        RECT 120.600 189.190 131.500 189.690 ;
        RECT 120.500 188.690 131.400 189.190 ;
        RECT 137.250 188.990 139.000 190.260 ;
        RECT 120.500 188.440 127.400 188.690 ;
        RECT 128.100 188.470 129.600 188.690 ;
        RECT 120.500 188.390 121.450 188.440 ;
        RECT 120.500 188.190 121.400 188.390 ;
        RECT 113.000 184.290 116.120 188.120 ;
        RECT 116.500 187.590 121.400 188.190 ;
        RECT 122.000 188.130 123.950 188.240 ;
        RECT 121.950 187.900 123.950 188.130 ;
        RECT 116.500 185.390 116.800 187.590 ;
        RECT 117.700 187.230 119.500 187.390 ;
        RECT 117.500 187.000 119.500 187.230 ;
        RECT 117.110 186.840 117.340 186.950 ;
        RECT 117.700 186.940 119.500 187.000 ;
        RECT 117.700 186.840 119.250 186.940 ;
        RECT 117.100 186.790 117.400 186.840 ;
        RECT 119.660 186.790 119.890 186.950 ;
        RECT 117.100 186.690 117.500 186.790 ;
        RECT 119.500 186.690 119.900 186.790 ;
        RECT 117.100 186.240 119.900 186.690 ;
        RECT 117.100 186.090 117.500 186.240 ;
        RECT 119.550 186.090 119.900 186.240 ;
        RECT 120.100 186.290 121.400 187.590 ;
        RECT 121.560 187.690 121.790 187.850 ;
        RECT 124.110 187.690 124.340 187.850 ;
        RECT 121.560 187.090 124.340 187.690 ;
        RECT 121.560 186.890 121.790 187.090 ;
        RECT 124.110 186.890 124.340 187.090 ;
        RECT 122.400 186.840 123.900 186.890 ;
        RECT 121.950 186.610 123.950 186.840 ;
        RECT 122.400 186.290 123.900 186.610 ;
        RECT 124.600 186.590 127.400 188.440 ;
        RECT 128.050 188.240 130.050 188.470 ;
        RECT 127.660 187.990 127.890 188.190 ;
        RECT 130.210 188.180 130.440 188.190 ;
        RECT 130.210 188.040 130.500 188.180 ;
        RECT 130.100 187.990 130.500 188.040 ;
        RECT 127.660 187.230 130.500 187.990 ;
        RECT 127.700 187.040 130.500 187.230 ;
        RECT 127.700 186.990 130.400 187.040 ;
        RECT 128.050 186.950 130.050 186.990 ;
        RECT 130.700 186.590 131.400 188.690 ;
        RECT 124.600 186.290 131.400 186.590 ;
        RECT 117.100 186.040 117.400 186.090 ;
        RECT 117.110 185.990 117.340 186.040 ;
        RECT 119.660 185.990 119.890 186.090 ;
        RECT 117.800 185.940 119.400 185.990 ;
        RECT 117.500 185.710 119.500 185.940 ;
        RECT 120.100 185.890 131.400 186.290 ;
        RECT 117.800 185.540 119.450 185.710 ;
        RECT 120.100 185.690 127.400 185.890 ;
        RECT 120.100 185.390 121.400 185.690 ;
        RECT 124.550 185.640 127.400 185.690 ;
        RECT 122.000 185.490 122.500 185.540 ;
        RECT 116.500 184.890 121.400 185.390 ;
        RECT 121.950 185.000 123.950 185.490 ;
        RECT 113.000 183.720 119.900 184.290 ;
        RECT 113.000 181.990 114.300 183.720 ;
        RECT 119.580 183.690 119.900 183.720 ;
        RECT 114.905 183.390 118.905 183.430 ;
        RECT 114.500 183.150 119.300 183.390 ;
        RECT 114.470 182.290 119.340 183.150 ;
        RECT 114.470 182.190 114.700 182.290 ;
        RECT 119.110 182.190 119.340 182.290 ;
        RECT 114.905 181.990 118.905 182.140 ;
        RECT 119.600 181.990 119.900 183.690 ;
        RECT 113.000 180.390 119.900 181.990 ;
        RECT 113.000 180.290 118.905 180.390 ;
        RECT 113.000 178.590 114.300 180.290 ;
        RECT 114.905 180.200 118.905 180.290 ;
        RECT 114.470 179.990 114.700 180.150 ;
        RECT 119.110 179.990 119.340 180.150 ;
        RECT 114.470 179.490 119.340 179.990 ;
        RECT 114.470 179.390 114.800 179.490 ;
        RECT 114.470 179.190 114.700 179.390 ;
        RECT 115.600 179.340 115.900 179.490 ;
        RECT 119.100 179.390 119.340 179.490 ;
        RECT 116.900 179.140 118.700 179.240 ;
        RECT 119.110 179.190 119.340 179.390 ;
        RECT 114.905 178.910 118.905 179.140 ;
        RECT 116.900 178.740 118.700 178.910 ;
        RECT 119.600 178.590 119.900 180.390 ;
        RECT 113.000 177.390 119.900 178.590 ;
        RECT 120.600 183.390 121.400 184.890 ;
        RECT 121.560 184.790 121.790 184.950 ;
        RECT 124.110 184.790 124.340 184.950 ;
        RECT 121.560 184.190 124.340 184.790 ;
        RECT 121.560 183.990 121.790 184.190 ;
        RECT 124.110 183.990 124.340 184.190 ;
        RECT 122.400 183.940 123.900 183.990 ;
        RECT 121.950 183.710 123.950 183.940 ;
        RECT 122.400 183.390 123.900 183.710 ;
        RECT 124.600 183.690 127.400 185.640 ;
        RECT 128.100 185.570 129.600 185.890 ;
        RECT 128.050 185.340 130.050 185.570 ;
        RECT 127.660 185.090 127.890 185.290 ;
        RECT 130.210 185.090 130.440 185.290 ;
        RECT 127.660 184.330 130.440 185.090 ;
        RECT 127.700 184.090 130.400 184.330 ;
        RECT 128.050 184.050 130.050 184.090 ;
        RECT 130.600 183.690 131.400 185.890 ;
        RECT 124.600 183.390 131.400 183.690 ;
        RECT 120.600 182.990 131.400 183.390 ;
        RECT 120.600 182.690 127.400 182.990 ;
        RECT 120.600 180.490 121.400 182.690 ;
        RECT 121.950 182.290 123.950 182.330 ;
        RECT 121.600 182.050 124.300 182.290 ;
        RECT 121.560 181.290 124.340 182.050 ;
        RECT 121.560 181.090 121.790 181.290 ;
        RECT 124.110 181.090 124.340 181.290 ;
        RECT 121.950 180.810 123.950 181.040 ;
        RECT 122.400 180.490 123.900 180.810 ;
        RECT 124.600 180.740 127.400 182.690 ;
        RECT 128.100 182.670 129.600 182.990 ;
        RECT 128.050 182.440 130.050 182.670 ;
        RECT 128.100 182.390 129.600 182.440 ;
        RECT 127.660 182.190 127.890 182.390 ;
        RECT 130.210 182.190 130.440 182.390 ;
        RECT 127.660 181.590 130.440 182.190 ;
        RECT 127.660 181.430 127.890 181.590 ;
        RECT 130.210 181.430 130.440 181.590 ;
        RECT 130.600 181.490 131.400 182.990 ;
        RECT 132.100 187.790 139.000 188.990 ;
        RECT 132.100 185.990 132.400 187.790 ;
        RECT 133.300 187.470 135.100 187.640 ;
        RECT 133.095 187.240 137.095 187.470 ;
        RECT 132.660 186.990 132.890 187.190 ;
        RECT 133.300 187.140 135.100 187.240 ;
        RECT 132.660 186.890 132.900 186.990 ;
        RECT 136.100 186.890 136.400 187.040 ;
        RECT 137.300 186.990 137.530 187.190 ;
        RECT 137.200 186.890 137.530 186.990 ;
        RECT 132.660 186.390 137.530 186.890 ;
        RECT 132.660 186.230 132.890 186.390 ;
        RECT 137.300 186.230 137.530 186.390 ;
        RECT 133.095 186.090 137.095 186.180 ;
        RECT 137.700 186.090 139.000 187.790 ;
        RECT 133.095 185.990 139.000 186.090 ;
        RECT 132.100 184.390 139.000 185.990 ;
        RECT 132.100 182.690 132.400 184.390 ;
        RECT 133.095 184.240 137.095 184.390 ;
        RECT 132.660 184.090 132.890 184.190 ;
        RECT 137.300 184.090 137.530 184.190 ;
        RECT 132.660 183.230 137.530 184.090 ;
        RECT 132.700 182.990 137.500 183.230 ;
        RECT 133.095 182.950 137.095 182.990 ;
        RECT 132.100 182.660 132.420 182.690 ;
        RECT 137.700 182.660 139.000 184.390 ;
        RECT 132.100 182.090 139.000 182.660 ;
        RECT 128.050 180.890 130.050 181.380 ;
        RECT 130.600 180.990 135.500 181.490 ;
        RECT 129.500 180.840 130.000 180.890 ;
        RECT 124.600 180.690 127.450 180.740 ;
        RECT 130.600 180.690 131.900 180.990 ;
        RECT 124.600 180.490 131.900 180.690 ;
        RECT 132.550 180.670 134.200 180.840 ;
        RECT 120.600 180.090 131.900 180.490 ;
        RECT 132.500 180.440 134.500 180.670 ;
        RECT 132.600 180.390 134.200 180.440 ;
        RECT 132.110 180.290 132.340 180.390 ;
        RECT 134.660 180.340 134.890 180.390 ;
        RECT 134.600 180.290 134.900 180.340 ;
        RECT 120.600 179.790 127.400 180.090 ;
        RECT 120.600 177.690 121.300 179.790 ;
        RECT 121.950 179.390 123.950 179.430 ;
        RECT 121.600 179.340 124.300 179.390 ;
        RECT 121.500 179.150 124.300 179.340 ;
        RECT 121.500 178.390 124.340 179.150 ;
        RECT 121.500 178.340 121.900 178.390 ;
        RECT 121.500 178.200 121.790 178.340 ;
        RECT 121.560 178.190 121.790 178.200 ;
        RECT 124.110 178.190 124.340 178.390 ;
        RECT 121.950 177.910 123.950 178.140 ;
        RECT 124.600 177.940 127.400 179.790 ;
        RECT 128.100 179.770 129.600 180.090 ;
        RECT 128.050 179.540 130.050 179.770 ;
        RECT 128.100 179.490 129.600 179.540 ;
        RECT 127.660 179.290 127.890 179.490 ;
        RECT 130.210 179.290 130.440 179.490 ;
        RECT 127.660 178.690 130.440 179.290 ;
        RECT 127.660 178.530 127.890 178.690 ;
        RECT 130.210 178.530 130.440 178.690 ;
        RECT 130.600 178.790 131.900 180.090 ;
        RECT 132.100 180.140 132.450 180.290 ;
        RECT 134.500 180.140 134.900 180.290 ;
        RECT 132.100 179.690 134.900 180.140 ;
        RECT 132.100 179.590 132.500 179.690 ;
        RECT 134.500 179.590 134.900 179.690 ;
        RECT 132.110 179.430 132.340 179.590 ;
        RECT 134.600 179.540 134.900 179.590 ;
        RECT 132.750 179.440 134.300 179.540 ;
        RECT 132.500 179.380 134.300 179.440 ;
        RECT 134.660 179.430 134.890 179.540 ;
        RECT 132.500 179.150 134.500 179.380 ;
        RECT 132.500 178.990 134.300 179.150 ;
        RECT 135.200 178.790 135.500 180.990 ;
        RECT 128.050 178.250 130.050 178.480 ;
        RECT 128.050 178.140 130.000 178.250 ;
        RECT 130.600 178.190 135.500 178.790 ;
        RECT 135.880 178.260 139.000 182.090 ;
        RECT 130.600 177.990 131.500 178.190 ;
        RECT 130.550 177.940 131.500 177.990 ;
        RECT 122.400 177.690 123.900 177.910 ;
        RECT 124.600 177.690 131.500 177.940 ;
        RECT 113.000 176.120 114.750 177.390 ;
        RECT 120.600 177.190 131.500 177.690 ;
        RECT 120.500 176.690 131.400 177.190 ;
        RECT 137.250 176.990 139.000 178.260 ;
        RECT 120.500 176.440 127.400 176.690 ;
        RECT 128.100 176.470 129.600 176.690 ;
        RECT 120.500 176.390 121.450 176.440 ;
        RECT 120.500 176.190 121.400 176.390 ;
        RECT 113.000 172.290 116.120 176.120 ;
        RECT 116.500 175.590 121.400 176.190 ;
        RECT 122.000 176.130 123.950 176.240 ;
        RECT 121.950 175.900 123.950 176.130 ;
        RECT 116.500 173.390 116.800 175.590 ;
        RECT 117.700 175.230 119.500 175.390 ;
        RECT 117.500 175.000 119.500 175.230 ;
        RECT 117.110 174.840 117.340 174.950 ;
        RECT 117.700 174.940 119.500 175.000 ;
        RECT 117.700 174.840 119.250 174.940 ;
        RECT 117.100 174.790 117.400 174.840 ;
        RECT 119.660 174.790 119.890 174.950 ;
        RECT 117.100 174.690 117.500 174.790 ;
        RECT 119.500 174.690 119.900 174.790 ;
        RECT 117.100 174.240 119.900 174.690 ;
        RECT 117.100 174.090 117.500 174.240 ;
        RECT 119.550 174.090 119.900 174.240 ;
        RECT 120.100 174.290 121.400 175.590 ;
        RECT 121.560 175.690 121.790 175.850 ;
        RECT 124.110 175.690 124.340 175.850 ;
        RECT 121.560 175.090 124.340 175.690 ;
        RECT 121.560 174.890 121.790 175.090 ;
        RECT 124.110 174.890 124.340 175.090 ;
        RECT 122.400 174.840 123.900 174.890 ;
        RECT 121.950 174.610 123.950 174.840 ;
        RECT 122.400 174.290 123.900 174.610 ;
        RECT 124.600 174.590 127.400 176.440 ;
        RECT 128.050 176.240 130.050 176.470 ;
        RECT 127.660 175.990 127.890 176.190 ;
        RECT 130.210 176.180 130.440 176.190 ;
        RECT 130.210 176.040 130.500 176.180 ;
        RECT 130.100 175.990 130.500 176.040 ;
        RECT 127.660 175.230 130.500 175.990 ;
        RECT 127.700 175.040 130.500 175.230 ;
        RECT 127.700 174.990 130.400 175.040 ;
        RECT 128.050 174.950 130.050 174.990 ;
        RECT 130.700 174.590 131.400 176.690 ;
        RECT 124.600 174.290 131.400 174.590 ;
        RECT 117.100 174.040 117.400 174.090 ;
        RECT 117.110 173.990 117.340 174.040 ;
        RECT 119.660 173.990 119.890 174.090 ;
        RECT 117.800 173.940 119.400 173.990 ;
        RECT 117.500 173.710 119.500 173.940 ;
        RECT 120.100 173.890 131.400 174.290 ;
        RECT 117.800 173.540 119.450 173.710 ;
        RECT 120.100 173.690 127.400 173.890 ;
        RECT 120.100 173.390 121.400 173.690 ;
        RECT 124.550 173.640 127.400 173.690 ;
        RECT 122.000 173.490 122.500 173.540 ;
        RECT 116.500 172.890 121.400 173.390 ;
        RECT 121.950 173.000 123.950 173.490 ;
        RECT 113.000 171.720 119.900 172.290 ;
        RECT 113.000 169.990 114.300 171.720 ;
        RECT 119.580 171.690 119.900 171.720 ;
        RECT 114.905 171.390 118.905 171.430 ;
        RECT 114.500 171.150 119.300 171.390 ;
        RECT 114.470 170.290 119.340 171.150 ;
        RECT 114.470 170.190 114.700 170.290 ;
        RECT 119.110 170.190 119.340 170.290 ;
        RECT 114.905 169.990 118.905 170.140 ;
        RECT 119.600 169.990 119.900 171.690 ;
        RECT 113.000 168.390 119.900 169.990 ;
        RECT 113.000 168.290 118.905 168.390 ;
        RECT 113.000 166.590 114.300 168.290 ;
        RECT 114.905 168.200 118.905 168.290 ;
        RECT 114.470 167.990 114.700 168.150 ;
        RECT 119.110 167.990 119.340 168.150 ;
        RECT 114.470 167.490 119.340 167.990 ;
        RECT 114.470 167.390 114.800 167.490 ;
        RECT 114.470 167.190 114.700 167.390 ;
        RECT 115.600 167.340 115.900 167.490 ;
        RECT 119.100 167.390 119.340 167.490 ;
        RECT 116.900 167.140 118.700 167.240 ;
        RECT 119.110 167.190 119.340 167.390 ;
        RECT 114.905 166.910 118.905 167.140 ;
        RECT 116.900 166.740 118.700 166.910 ;
        RECT 119.600 166.590 119.900 168.390 ;
        RECT 113.000 165.390 119.900 166.590 ;
        RECT 120.600 171.390 121.400 172.890 ;
        RECT 121.560 172.790 121.790 172.950 ;
        RECT 124.110 172.790 124.340 172.950 ;
        RECT 121.560 172.190 124.340 172.790 ;
        RECT 121.560 171.990 121.790 172.190 ;
        RECT 124.110 171.990 124.340 172.190 ;
        RECT 122.400 171.940 123.900 171.990 ;
        RECT 121.950 171.710 123.950 171.940 ;
        RECT 122.400 171.390 123.900 171.710 ;
        RECT 124.600 171.690 127.400 173.640 ;
        RECT 128.100 173.570 129.600 173.890 ;
        RECT 128.050 173.340 130.050 173.570 ;
        RECT 127.660 173.090 127.890 173.290 ;
        RECT 130.210 173.090 130.440 173.290 ;
        RECT 127.660 172.330 130.440 173.090 ;
        RECT 127.700 172.090 130.400 172.330 ;
        RECT 128.050 172.050 130.050 172.090 ;
        RECT 130.600 171.690 131.400 173.890 ;
        RECT 124.600 171.390 131.400 171.690 ;
        RECT 120.600 170.990 131.400 171.390 ;
        RECT 120.600 170.690 127.400 170.990 ;
        RECT 120.600 168.490 121.400 170.690 ;
        RECT 121.950 170.290 123.950 170.330 ;
        RECT 121.600 170.050 124.300 170.290 ;
        RECT 121.560 169.290 124.340 170.050 ;
        RECT 121.560 169.090 121.790 169.290 ;
        RECT 124.110 169.090 124.340 169.290 ;
        RECT 121.950 168.810 123.950 169.040 ;
        RECT 122.400 168.490 123.900 168.810 ;
        RECT 124.600 168.740 127.400 170.690 ;
        RECT 128.100 170.670 129.600 170.990 ;
        RECT 128.050 170.440 130.050 170.670 ;
        RECT 128.100 170.390 129.600 170.440 ;
        RECT 127.660 170.190 127.890 170.390 ;
        RECT 130.210 170.190 130.440 170.390 ;
        RECT 127.660 169.590 130.440 170.190 ;
        RECT 127.660 169.430 127.890 169.590 ;
        RECT 130.210 169.430 130.440 169.590 ;
        RECT 130.600 169.490 131.400 170.990 ;
        RECT 132.100 175.790 139.000 176.990 ;
        RECT 132.100 173.990 132.400 175.790 ;
        RECT 133.300 175.470 135.100 175.640 ;
        RECT 133.095 175.240 137.095 175.470 ;
        RECT 132.660 174.990 132.890 175.190 ;
        RECT 133.300 175.140 135.100 175.240 ;
        RECT 132.660 174.890 132.900 174.990 ;
        RECT 136.100 174.890 136.400 175.040 ;
        RECT 137.300 174.990 137.530 175.190 ;
        RECT 137.200 174.890 137.530 174.990 ;
        RECT 132.660 174.390 137.530 174.890 ;
        RECT 132.660 174.230 132.890 174.390 ;
        RECT 137.300 174.230 137.530 174.390 ;
        RECT 133.095 174.090 137.095 174.180 ;
        RECT 137.700 174.090 139.000 175.790 ;
        RECT 133.095 173.990 139.000 174.090 ;
        RECT 132.100 172.390 139.000 173.990 ;
        RECT 132.100 170.690 132.400 172.390 ;
        RECT 133.095 172.240 137.095 172.390 ;
        RECT 132.660 172.090 132.890 172.190 ;
        RECT 137.300 172.090 137.530 172.190 ;
        RECT 132.660 171.230 137.530 172.090 ;
        RECT 132.700 170.990 137.500 171.230 ;
        RECT 133.095 170.950 137.095 170.990 ;
        RECT 132.100 170.660 132.420 170.690 ;
        RECT 137.700 170.660 139.000 172.390 ;
        RECT 132.100 170.090 139.000 170.660 ;
        RECT 128.050 168.890 130.050 169.380 ;
        RECT 130.600 168.990 135.500 169.490 ;
        RECT 129.500 168.840 130.000 168.890 ;
        RECT 124.600 168.690 127.450 168.740 ;
        RECT 130.600 168.690 131.900 168.990 ;
        RECT 124.600 168.490 131.900 168.690 ;
        RECT 132.550 168.670 134.200 168.840 ;
        RECT 120.600 168.090 131.900 168.490 ;
        RECT 132.500 168.440 134.500 168.670 ;
        RECT 132.600 168.390 134.200 168.440 ;
        RECT 132.110 168.290 132.340 168.390 ;
        RECT 134.660 168.340 134.890 168.390 ;
        RECT 134.600 168.290 134.900 168.340 ;
        RECT 120.600 167.790 127.400 168.090 ;
        RECT 120.600 165.690 121.300 167.790 ;
        RECT 121.950 167.390 123.950 167.430 ;
        RECT 121.600 167.340 124.300 167.390 ;
        RECT 121.500 167.150 124.300 167.340 ;
        RECT 121.500 166.390 124.340 167.150 ;
        RECT 121.500 166.340 121.900 166.390 ;
        RECT 121.500 166.200 121.790 166.340 ;
        RECT 121.560 166.190 121.790 166.200 ;
        RECT 124.110 166.190 124.340 166.390 ;
        RECT 121.950 165.910 123.950 166.140 ;
        RECT 124.600 165.940 127.400 167.790 ;
        RECT 128.100 167.770 129.600 168.090 ;
        RECT 128.050 167.540 130.050 167.770 ;
        RECT 128.100 167.490 129.600 167.540 ;
        RECT 127.660 167.290 127.890 167.490 ;
        RECT 130.210 167.290 130.440 167.490 ;
        RECT 127.660 166.690 130.440 167.290 ;
        RECT 127.660 166.530 127.890 166.690 ;
        RECT 130.210 166.530 130.440 166.690 ;
        RECT 130.600 166.790 131.900 168.090 ;
        RECT 132.100 168.140 132.450 168.290 ;
        RECT 134.500 168.140 134.900 168.290 ;
        RECT 132.100 167.690 134.900 168.140 ;
        RECT 132.100 167.590 132.500 167.690 ;
        RECT 134.500 167.590 134.900 167.690 ;
        RECT 132.110 167.430 132.340 167.590 ;
        RECT 134.600 167.540 134.900 167.590 ;
        RECT 132.750 167.440 134.300 167.540 ;
        RECT 132.500 167.380 134.300 167.440 ;
        RECT 134.660 167.430 134.890 167.540 ;
        RECT 132.500 167.150 134.500 167.380 ;
        RECT 132.500 166.990 134.300 167.150 ;
        RECT 135.200 166.790 135.500 168.990 ;
        RECT 128.050 166.250 130.050 166.480 ;
        RECT 128.050 166.140 130.000 166.250 ;
        RECT 130.600 166.190 135.500 166.790 ;
        RECT 135.880 166.260 139.000 170.090 ;
        RECT 130.600 165.990 131.500 166.190 ;
        RECT 130.550 165.940 131.500 165.990 ;
        RECT 122.400 165.690 123.900 165.910 ;
        RECT 124.600 165.690 131.500 165.940 ;
        RECT 113.000 164.120 114.750 165.390 ;
        RECT 120.600 165.190 131.500 165.690 ;
        RECT 120.500 164.690 131.400 165.190 ;
        RECT 137.250 164.990 139.000 166.260 ;
        RECT 120.500 164.440 127.400 164.690 ;
        RECT 128.100 164.470 129.600 164.690 ;
        RECT 120.500 164.390 121.450 164.440 ;
        RECT 120.500 164.190 121.400 164.390 ;
        RECT 113.000 160.290 116.120 164.120 ;
        RECT 116.500 163.590 121.400 164.190 ;
        RECT 122.000 164.130 123.950 164.240 ;
        RECT 121.950 163.900 123.950 164.130 ;
        RECT 116.500 161.390 116.800 163.590 ;
        RECT 117.700 163.230 119.500 163.390 ;
        RECT 117.500 163.000 119.500 163.230 ;
        RECT 117.110 162.840 117.340 162.950 ;
        RECT 117.700 162.940 119.500 163.000 ;
        RECT 117.700 162.840 119.250 162.940 ;
        RECT 117.100 162.790 117.400 162.840 ;
        RECT 119.660 162.790 119.890 162.950 ;
        RECT 117.100 162.690 117.500 162.790 ;
        RECT 119.500 162.690 119.900 162.790 ;
        RECT 117.100 162.240 119.900 162.690 ;
        RECT 117.100 162.090 117.500 162.240 ;
        RECT 119.550 162.090 119.900 162.240 ;
        RECT 120.100 162.290 121.400 163.590 ;
        RECT 121.560 163.690 121.790 163.850 ;
        RECT 124.110 163.690 124.340 163.850 ;
        RECT 121.560 163.090 124.340 163.690 ;
        RECT 121.560 162.890 121.790 163.090 ;
        RECT 124.110 162.890 124.340 163.090 ;
        RECT 122.400 162.840 123.900 162.890 ;
        RECT 121.950 162.610 123.950 162.840 ;
        RECT 122.400 162.290 123.900 162.610 ;
        RECT 124.600 162.590 127.400 164.440 ;
        RECT 128.050 164.240 130.050 164.470 ;
        RECT 127.660 163.990 127.890 164.190 ;
        RECT 130.210 164.180 130.440 164.190 ;
        RECT 130.210 164.040 130.500 164.180 ;
        RECT 130.100 163.990 130.500 164.040 ;
        RECT 127.660 163.230 130.500 163.990 ;
        RECT 127.700 163.040 130.500 163.230 ;
        RECT 127.700 162.990 130.400 163.040 ;
        RECT 128.050 162.950 130.050 162.990 ;
        RECT 130.700 162.590 131.400 164.690 ;
        RECT 124.600 162.290 131.400 162.590 ;
        RECT 117.100 162.040 117.400 162.090 ;
        RECT 117.110 161.990 117.340 162.040 ;
        RECT 119.660 161.990 119.890 162.090 ;
        RECT 117.800 161.940 119.400 161.990 ;
        RECT 117.500 161.710 119.500 161.940 ;
        RECT 120.100 161.890 131.400 162.290 ;
        RECT 117.800 161.540 119.450 161.710 ;
        RECT 120.100 161.690 127.400 161.890 ;
        RECT 120.100 161.390 121.400 161.690 ;
        RECT 124.550 161.640 127.400 161.690 ;
        RECT 122.000 161.490 122.500 161.540 ;
        RECT 116.500 160.890 121.400 161.390 ;
        RECT 121.950 161.000 123.950 161.490 ;
        RECT 113.000 159.720 119.900 160.290 ;
        RECT 113.000 157.990 114.300 159.720 ;
        RECT 119.580 159.690 119.900 159.720 ;
        RECT 114.905 159.390 118.905 159.430 ;
        RECT 114.500 159.150 119.300 159.390 ;
        RECT 114.470 158.290 119.340 159.150 ;
        RECT 114.470 158.190 114.700 158.290 ;
        RECT 119.110 158.190 119.340 158.290 ;
        RECT 114.905 157.990 118.905 158.140 ;
        RECT 119.600 157.990 119.900 159.690 ;
        RECT 113.000 156.390 119.900 157.990 ;
        RECT 113.000 156.290 118.905 156.390 ;
        RECT 113.000 154.590 114.300 156.290 ;
        RECT 114.905 156.200 118.905 156.290 ;
        RECT 114.470 155.990 114.700 156.150 ;
        RECT 119.110 155.990 119.340 156.150 ;
        RECT 114.470 155.490 119.340 155.990 ;
        RECT 114.470 155.390 114.800 155.490 ;
        RECT 114.470 155.190 114.700 155.390 ;
        RECT 115.600 155.340 115.900 155.490 ;
        RECT 119.100 155.390 119.340 155.490 ;
        RECT 116.900 155.140 118.700 155.240 ;
        RECT 119.110 155.190 119.340 155.390 ;
        RECT 114.905 154.910 118.905 155.140 ;
        RECT 116.900 154.740 118.700 154.910 ;
        RECT 119.600 154.590 119.900 156.390 ;
        RECT 113.000 153.390 119.900 154.590 ;
        RECT 120.600 159.390 121.400 160.890 ;
        RECT 121.560 160.790 121.790 160.950 ;
        RECT 124.110 160.790 124.340 160.950 ;
        RECT 121.560 160.190 124.340 160.790 ;
        RECT 121.560 159.990 121.790 160.190 ;
        RECT 124.110 159.990 124.340 160.190 ;
        RECT 122.400 159.940 123.900 159.990 ;
        RECT 121.950 159.710 123.950 159.940 ;
        RECT 122.400 159.390 123.900 159.710 ;
        RECT 124.600 159.690 127.400 161.640 ;
        RECT 128.100 161.570 129.600 161.890 ;
        RECT 128.050 161.340 130.050 161.570 ;
        RECT 127.660 161.090 127.890 161.290 ;
        RECT 130.210 161.090 130.440 161.290 ;
        RECT 127.660 160.330 130.440 161.090 ;
        RECT 127.700 160.090 130.400 160.330 ;
        RECT 128.050 160.050 130.050 160.090 ;
        RECT 130.600 159.690 131.400 161.890 ;
        RECT 124.600 159.390 131.400 159.690 ;
        RECT 120.600 158.990 131.400 159.390 ;
        RECT 120.600 158.690 127.400 158.990 ;
        RECT 120.600 156.490 121.400 158.690 ;
        RECT 121.950 158.290 123.950 158.330 ;
        RECT 121.600 158.050 124.300 158.290 ;
        RECT 121.560 157.290 124.340 158.050 ;
        RECT 121.560 157.090 121.790 157.290 ;
        RECT 124.110 157.090 124.340 157.290 ;
        RECT 121.950 156.810 123.950 157.040 ;
        RECT 122.400 156.490 123.900 156.810 ;
        RECT 124.600 156.740 127.400 158.690 ;
        RECT 128.100 158.670 129.600 158.990 ;
        RECT 128.050 158.440 130.050 158.670 ;
        RECT 128.100 158.390 129.600 158.440 ;
        RECT 127.660 158.190 127.890 158.390 ;
        RECT 130.210 158.190 130.440 158.390 ;
        RECT 127.660 157.590 130.440 158.190 ;
        RECT 127.660 157.430 127.890 157.590 ;
        RECT 130.210 157.430 130.440 157.590 ;
        RECT 130.600 157.490 131.400 158.990 ;
        RECT 132.100 163.790 139.000 164.990 ;
        RECT 132.100 161.990 132.400 163.790 ;
        RECT 133.300 163.470 135.100 163.640 ;
        RECT 133.095 163.240 137.095 163.470 ;
        RECT 132.660 162.990 132.890 163.190 ;
        RECT 133.300 163.140 135.100 163.240 ;
        RECT 132.660 162.890 132.900 162.990 ;
        RECT 136.100 162.890 136.400 163.040 ;
        RECT 137.300 162.990 137.530 163.190 ;
        RECT 137.200 162.890 137.530 162.990 ;
        RECT 132.660 162.390 137.530 162.890 ;
        RECT 132.660 162.230 132.890 162.390 ;
        RECT 137.300 162.230 137.530 162.390 ;
        RECT 133.095 162.090 137.095 162.180 ;
        RECT 137.700 162.090 139.000 163.790 ;
        RECT 133.095 161.990 139.000 162.090 ;
        RECT 132.100 160.390 139.000 161.990 ;
        RECT 132.100 158.690 132.400 160.390 ;
        RECT 133.095 160.240 137.095 160.390 ;
        RECT 132.660 160.090 132.890 160.190 ;
        RECT 137.300 160.090 137.530 160.190 ;
        RECT 132.660 159.230 137.530 160.090 ;
        RECT 132.700 158.990 137.500 159.230 ;
        RECT 133.095 158.950 137.095 158.990 ;
        RECT 132.100 158.660 132.420 158.690 ;
        RECT 137.700 158.660 139.000 160.390 ;
        RECT 132.100 158.090 139.000 158.660 ;
        RECT 128.050 156.890 130.050 157.380 ;
        RECT 130.600 156.990 135.500 157.490 ;
        RECT 129.500 156.840 130.000 156.890 ;
        RECT 124.600 156.690 127.450 156.740 ;
        RECT 130.600 156.690 131.900 156.990 ;
        RECT 124.600 156.490 131.900 156.690 ;
        RECT 132.550 156.670 134.200 156.840 ;
        RECT 120.600 156.090 131.900 156.490 ;
        RECT 132.500 156.440 134.500 156.670 ;
        RECT 132.600 156.390 134.200 156.440 ;
        RECT 132.110 156.290 132.340 156.390 ;
        RECT 134.660 156.340 134.890 156.390 ;
        RECT 134.600 156.290 134.900 156.340 ;
        RECT 120.600 155.790 127.400 156.090 ;
        RECT 120.600 153.690 121.300 155.790 ;
        RECT 121.950 155.390 123.950 155.430 ;
        RECT 121.600 155.340 124.300 155.390 ;
        RECT 121.500 155.150 124.300 155.340 ;
        RECT 121.500 154.390 124.340 155.150 ;
        RECT 121.500 154.340 121.900 154.390 ;
        RECT 121.500 154.200 121.790 154.340 ;
        RECT 121.560 154.190 121.790 154.200 ;
        RECT 124.110 154.190 124.340 154.390 ;
        RECT 121.950 153.910 123.950 154.140 ;
        RECT 124.600 153.940 127.400 155.790 ;
        RECT 128.100 155.770 129.600 156.090 ;
        RECT 128.050 155.540 130.050 155.770 ;
        RECT 128.100 155.490 129.600 155.540 ;
        RECT 127.660 155.290 127.890 155.490 ;
        RECT 130.210 155.290 130.440 155.490 ;
        RECT 127.660 154.690 130.440 155.290 ;
        RECT 127.660 154.530 127.890 154.690 ;
        RECT 130.210 154.530 130.440 154.690 ;
        RECT 130.600 154.790 131.900 156.090 ;
        RECT 132.100 156.140 132.450 156.290 ;
        RECT 134.500 156.140 134.900 156.290 ;
        RECT 132.100 155.690 134.900 156.140 ;
        RECT 132.100 155.590 132.500 155.690 ;
        RECT 134.500 155.590 134.900 155.690 ;
        RECT 132.110 155.430 132.340 155.590 ;
        RECT 134.600 155.540 134.900 155.590 ;
        RECT 132.750 155.440 134.300 155.540 ;
        RECT 132.500 155.380 134.300 155.440 ;
        RECT 134.660 155.430 134.890 155.540 ;
        RECT 132.500 155.150 134.500 155.380 ;
        RECT 132.500 154.990 134.300 155.150 ;
        RECT 135.200 154.790 135.500 156.990 ;
        RECT 128.050 154.250 130.050 154.480 ;
        RECT 128.050 154.140 130.000 154.250 ;
        RECT 130.600 154.190 135.500 154.790 ;
        RECT 135.880 154.260 139.000 158.090 ;
        RECT 130.600 153.990 131.500 154.190 ;
        RECT 130.550 153.940 131.500 153.990 ;
        RECT 122.400 153.690 123.900 153.910 ;
        RECT 124.600 153.690 131.500 153.940 ;
        RECT 113.000 153.190 114.750 153.390 ;
        RECT 120.600 153.190 131.500 153.690 ;
        RECT 137.250 153.190 139.000 154.260 ;
        RECT 113.000 152.190 114.500 153.190 ;
        RECT 120.500 152.690 131.500 153.190 ;
        RECT 137.255 152.690 139.000 153.190 ;
        RECT 139.500 152.690 142.500 203.890 ;
        RECT 113.000 151.790 119.500 152.190 ;
        RECT 110.100 151.690 119.500 151.790 ;
        RECT 120.500 151.690 135.300 152.690 ;
        RECT 110.100 151.290 119.900 151.690 ;
        RECT 110.100 151.090 131.700 151.290 ;
        RECT 110.100 150.890 131.800 151.090 ;
        RECT 110.100 150.490 120.400 150.890 ;
        RECT 120.850 150.820 131.800 150.890 ;
        RECT 123.500 150.790 131.800 150.820 ;
        RECT 110.100 149.690 120.300 150.490 ;
        RECT 121.100 150.480 125.000 150.490 ;
        RECT 121.100 150.250 125.105 150.480 ;
        RECT 110.000 149.090 120.300 149.690 ;
        RECT 120.670 149.890 120.900 150.200 ;
        RECT 121.100 149.890 125.000 150.250 ;
        RECT 125.310 150.090 125.540 150.200 ;
        RECT 126.220 150.090 126.450 150.200 ;
        RECT 125.310 149.890 126.450 150.090 ;
        RECT 126.600 150.040 130.700 150.590 ;
        RECT 130.860 149.890 131.090 150.200 ;
        RECT 120.670 149.490 131.090 149.890 ;
        RECT 120.670 149.240 120.900 149.490 ;
        RECT 125.310 149.390 131.090 149.490 ;
        RECT 125.310 149.290 126.450 149.390 ;
        RECT 125.310 149.240 125.540 149.290 ;
        RECT 126.220 149.240 126.450 149.290 ;
        RECT 130.860 149.240 131.090 149.390 ;
        RECT 110.000 148.690 120.400 149.090 ;
        RECT 121.105 148.960 125.105 149.190 ;
        RECT 126.655 148.960 130.655 149.190 ;
        RECT 121.600 148.690 124.700 148.960 ;
        RECT 126.800 148.690 130.500 148.960 ;
        RECT 131.300 148.690 131.800 150.790 ;
        RECT 132.400 149.490 135.300 151.690 ;
        RECT 137.255 151.190 142.500 152.690 ;
        RECT 137.500 148.690 142.500 151.190 ;
        RECT 110.000 146.890 142.500 148.690 ;
        RECT 110.000 146.190 126.400 146.890 ;
        RECT 130.300 146.190 142.500 146.890 ;
        RECT 113.000 131.350 113.960 131.530 ;
        RECT 113.000 131.300 114.250 131.350 ;
        RECT 112.720 130.100 112.950 131.095 ;
        RECT 112.000 129.650 112.950 130.100 ;
        RECT 111.120 128.850 112.950 129.650 ;
        RECT 112.000 128.700 112.950 128.850 ;
        RECT 112.720 127.095 112.950 128.700 ;
        RECT 113.100 126.890 114.250 131.300 ;
        RECT 113.000 126.700 114.250 126.890 ;
        RECT 113.000 126.660 113.960 126.700 ;
        RECT 105.050 62.950 143.050 67.000 ;
        RECT 105.050 61.700 118.050 62.950 ;
        RECT 118.950 62.530 121.250 62.600 ;
        RECT 118.950 62.300 121.300 62.530 ;
        RECT 118.770 61.700 119.000 62.095 ;
        RECT 105.050 51.500 119.000 61.700 ;
        RECT 108.050 51.400 119.000 51.500 ;
        RECT 105.050 48.500 106.050 51.000 ;
        RECT 106.550 50.500 107.550 51.000 ;
        RECT 106.500 49.500 107.600 50.500 ;
        RECT 105.000 47.500 106.100 48.500 ;
        RECT 105.050 40.500 106.050 47.500 ;
        RECT 106.550 42.000 107.550 49.500 ;
        RECT 108.050 45.400 108.550 51.400 ;
        RECT 111.150 51.000 119.000 51.400 ;
        RECT 109.150 50.780 109.750 50.800 ;
        RECT 109.150 50.550 110.420 50.780 ;
        RECT 109.150 46.140 109.750 50.550 ;
        RECT 110.470 49.850 110.700 50.345 ;
        RECT 111.150 49.850 113.050 51.000 ;
        RECT 114.050 50.700 115.010 50.710 ;
        RECT 113.750 50.480 115.010 50.700 ;
        RECT 113.750 49.850 114.350 50.480 ;
        RECT 115.060 50.200 115.290 50.275 ;
        RECT 110.470 46.700 114.350 49.850 ;
        RECT 114.900 49.500 115.400 50.200 ;
        RECT 110.470 46.345 110.700 46.700 ;
        RECT 109.150 45.910 110.420 46.140 ;
        RECT 109.150 45.900 109.750 45.910 ;
        RECT 111.150 45.400 113.050 46.700 ;
        RECT 113.750 46.070 114.350 46.700 ;
        RECT 115.060 46.275 115.290 49.500 ;
        RECT 116.050 46.250 119.000 51.000 ;
        RECT 119.350 50.500 119.550 62.300 ;
        RECT 120.060 61.800 120.290 62.095 ;
        RECT 119.750 50.900 120.550 61.800 ;
        RECT 119.250 48.500 119.750 50.500 ;
        RECT 119.200 47.500 119.800 48.500 ;
        RECT 113.750 45.840 115.010 46.070 ;
        RECT 113.750 45.800 114.350 45.840 ;
        RECT 116.050 45.400 118.050 46.250 ;
        RECT 118.770 46.095 119.000 46.250 ;
        RECT 119.250 45.900 119.750 47.500 ;
        RECT 120.060 46.095 120.290 50.900 ;
        RECT 120.850 50.500 121.050 62.300 ;
        RECT 120.550 48.500 121.050 50.500 ;
        RECT 120.500 47.500 121.050 48.500 ;
        RECT 120.550 45.900 121.050 47.500 ;
        RECT 121.350 61.850 121.580 62.095 ;
        RECT 121.950 61.850 124.450 62.950 ;
        RECT 125.050 62.300 127.350 62.600 ;
        RECT 124.770 61.850 125.000 62.095 ;
        RECT 121.350 52.200 125.000 61.850 ;
        RECT 121.350 51.400 122.250 52.200 ;
        RECT 121.350 46.450 122.150 51.400 ;
        RECT 122.600 50.800 123.700 51.700 ;
        RECT 124.050 51.400 125.000 52.200 ;
        RECT 121.350 46.095 121.580 46.450 ;
        RECT 119.150 45.890 121.250 45.900 ;
        RECT 119.050 45.660 121.300 45.890 ;
        RECT 119.150 45.500 121.250 45.660 ;
        RECT 108.050 45.300 118.050 45.400 ;
        RECT 121.950 45.300 122.150 46.450 ;
        RECT 108.050 45.000 122.150 45.300 ;
        RECT 122.650 44.800 123.650 50.800 ;
        RECT 124.150 46.450 125.000 51.400 ;
        RECT 125.350 50.500 125.550 62.300 ;
        RECT 126.060 61.700 126.290 62.095 ;
        RECT 125.750 50.800 126.550 61.700 ;
        RECT 125.300 49.500 125.850 50.500 ;
        RECT 124.150 45.300 124.450 46.450 ;
        RECT 124.770 46.095 125.000 46.450 ;
        RECT 125.350 45.900 125.850 49.500 ;
        RECT 126.060 46.095 126.290 50.800 ;
        RECT 126.850 50.500 127.050 62.300 ;
        RECT 127.550 62.095 130.350 62.950 ;
        RECT 131.050 62.300 133.350 62.600 ;
        RECT 126.500 49.500 127.050 50.500 ;
        RECT 126.550 45.900 127.050 49.500 ;
        RECT 127.350 61.800 130.350 62.095 ;
        RECT 130.770 61.800 131.000 62.095 ;
        RECT 127.350 52.500 131.000 61.800 ;
        RECT 127.350 46.095 128.450 52.500 ;
        RECT 128.750 51.700 129.750 52.100 ;
        RECT 128.700 50.800 129.800 51.700 ;
        RECT 125.150 45.890 127.250 45.900 ;
        RECT 125.050 45.660 127.300 45.890 ;
        RECT 125.150 45.500 127.250 45.660 ;
        RECT 127.550 45.300 128.450 46.095 ;
        RECT 124.150 45.000 128.450 45.300 ;
        RECT 122.600 43.800 127.500 44.800 ;
        RECT 128.750 44.700 129.750 50.800 ;
        RECT 130.050 46.550 131.000 52.500 ;
        RECT 131.350 50.500 131.550 62.300 ;
        RECT 132.060 61.800 132.290 62.095 ;
        RECT 131.850 50.900 132.650 61.800 ;
        RECT 131.300 49.500 131.850 50.500 ;
        RECT 130.050 45.300 130.350 46.550 ;
        RECT 130.770 46.095 131.000 46.550 ;
        RECT 131.350 45.900 131.850 49.500 ;
        RECT 132.060 46.095 132.290 50.900 ;
        RECT 132.850 50.500 133.050 62.300 ;
        RECT 132.500 49.500 133.050 50.500 ;
        RECT 132.550 45.900 133.050 49.500 ;
        RECT 133.350 61.450 133.580 62.095 ;
        RECT 134.350 61.450 143.050 62.950 ;
        RECT 133.350 46.400 143.050 61.450 ;
        RECT 133.350 46.095 133.580 46.400 ;
        RECT 131.150 45.890 133.250 45.900 ;
        RECT 131.050 45.660 133.300 45.890 ;
        RECT 131.150 45.500 133.250 45.660 ;
        RECT 135.050 45.300 137.000 46.400 ;
        RECT 130.050 45.000 137.000 45.300 ;
        RECT 128.700 43.700 132.850 44.700 ;
        RECT 108.050 42.700 137.050 43.200 ;
        RECT 108.050 42.500 108.650 42.700 ;
        RECT 110.450 42.500 112.250 42.700 ;
        RECT 114.620 42.500 117.350 42.700 ;
        RECT 119.750 42.500 121.350 42.700 ;
        RECT 106.500 41.000 107.600 42.000 ;
        RECT 105.000 39.500 106.100 40.500 ;
        RECT 106.550 39.500 107.550 41.000 ;
        RECT 108.050 39.000 108.430 42.500 ;
        RECT 109.050 42.210 110.010 42.440 ;
        RECT 105.050 33.600 108.430 39.000 ;
        RECT 108.770 40.200 109.000 42.050 ;
        RECT 109.150 40.700 109.850 42.210 ;
        RECT 108.770 39.600 109.300 40.200 ;
        RECT 108.770 34.050 109.000 39.600 ;
        RECT 109.450 39.400 109.850 40.700 ;
        RECT 109.150 33.890 109.850 39.400 ;
        RECT 110.060 35.600 110.290 42.050 ;
        RECT 110.000 35.200 110.500 35.600 ;
        RECT 110.060 34.050 110.290 35.200 ;
        RECT 109.050 33.660 110.010 33.890 ;
        RECT 110.700 33.600 112.430 42.500 ;
        RECT 113.050 42.210 114.010 42.440 ;
        RECT 112.770 35.600 113.000 42.050 ;
        RECT 113.200 42.000 113.900 42.210 ;
        RECT 113.200 41.000 113.750 42.000 ;
        RECT 114.060 41.900 114.290 42.050 ;
        RECT 114.000 41.100 114.400 41.900 ;
        RECT 113.200 35.900 113.900 41.000 ;
        RECT 112.700 35.200 113.200 35.600 ;
        RECT 112.770 34.050 113.000 35.200 ;
        RECT 113.350 34.900 113.900 35.900 ;
        RECT 113.200 33.890 113.900 34.900 ;
        RECT 114.060 34.050 114.290 41.100 ;
        RECT 113.050 33.660 114.010 33.890 ;
        RECT 114.620 33.840 117.430 42.500 ;
        RECT 118.050 42.210 119.010 42.440 ;
        RECT 117.770 40.500 118.000 42.050 ;
        RECT 118.200 40.700 118.900 42.210 ;
        RECT 117.700 39.500 118.100 40.500 ;
        RECT 117.770 34.050 118.000 39.500 ;
        RECT 118.350 39.300 118.900 40.700 ;
        RECT 118.200 36.000 118.900 39.300 ;
        RECT 118.200 34.800 118.650 36.000 ;
        RECT 119.060 35.500 119.290 42.050 ;
        RECT 118.850 35.100 119.300 35.500 ;
        RECT 118.200 33.890 118.900 34.800 ;
        RECT 119.060 34.050 119.290 35.100 ;
        RECT 114.650 33.600 117.430 33.840 ;
        RECT 118.050 33.660 119.010 33.890 ;
        RECT 119.630 33.600 121.430 42.500 ;
        RECT 122.200 42.440 122.900 42.450 ;
        RECT 122.050 42.210 123.010 42.440 ;
        RECT 121.770 35.500 122.000 42.050 ;
        RECT 122.200 42.000 122.900 42.210 ;
        RECT 122.200 40.900 122.850 42.000 ;
        RECT 123.060 41.900 123.290 42.050 ;
        RECT 123.000 41.000 123.400 41.900 ;
        RECT 122.200 36.200 122.900 40.900 ;
        RECT 121.770 35.100 122.300 35.500 ;
        RECT 121.770 34.050 122.000 35.100 ;
        RECT 122.450 34.700 122.900 36.200 ;
        RECT 122.200 33.890 122.900 34.700 ;
        RECT 123.060 34.050 123.290 41.000 ;
        RECT 122.050 33.660 123.010 33.890 ;
        RECT 105.050 33.300 108.350 33.600 ;
        RECT 110.700 33.300 112.250 33.600 ;
        RECT 114.650 33.300 117.250 33.600 ;
        RECT 119.850 33.300 121.350 33.600 ;
        RECT 123.650 33.300 126.350 42.700 ;
        RECT 127.050 42.210 128.010 42.440 ;
        RECT 126.770 41.200 127.000 42.050 ;
        RECT 128.060 41.600 128.290 42.050 ;
        RECT 129.050 41.600 130.050 42.700 ;
        RECT 131.350 42.440 133.050 42.500 ;
        RECT 131.050 42.210 133.300 42.440 ;
        RECT 131.250 42.200 133.050 42.210 ;
        RECT 130.770 41.600 131.000 42.050 ;
        RECT 105.050 30.900 126.350 33.300 ;
        RECT 105.050 13.550 108.250 30.900 ;
        RECT 114.300 30.650 126.350 30.900 ;
        RECT 108.870 30.400 109.830 30.630 ;
        RECT 110.160 30.400 111.120 30.630 ;
        RECT 111.450 30.400 112.410 30.630 ;
        RECT 112.740 30.400 113.700 30.630 ;
        RECT 108.590 27.700 108.820 30.240 ;
        RECT 109.100 27.800 109.520 30.400 ;
        RECT 108.550 26.500 109.000 27.700 ;
        RECT 108.590 14.240 108.820 26.500 ;
        RECT 109.200 26.250 109.520 27.800 ;
        RECT 109.100 14.080 109.520 26.250 ;
        RECT 109.880 16.250 110.110 30.240 ;
        RECT 110.450 28.100 110.870 30.400 ;
        RECT 110.450 28.000 110.750 28.100 ;
        RECT 110.250 26.100 110.750 28.000 ;
        RECT 111.170 27.400 111.400 30.240 ;
        RECT 111.650 27.800 112.070 30.400 ;
        RECT 111.650 27.600 112.150 27.800 ;
        RECT 111.000 26.700 111.600 27.400 ;
        RECT 110.250 26.000 110.870 26.100 ;
        RECT 110.450 22.500 110.870 26.000 ;
        RECT 110.450 21.900 110.900 22.500 ;
        RECT 109.700 15.500 110.300 16.250 ;
        RECT 109.880 14.240 110.110 15.500 ;
        RECT 110.450 14.080 110.870 21.900 ;
        RECT 111.170 14.240 111.400 26.700 ;
        RECT 111.750 26.500 112.150 27.600 ;
        RECT 111.650 26.400 112.150 26.500 ;
        RECT 111.650 22.600 112.070 26.400 ;
        RECT 111.650 22.000 112.100 22.600 ;
        RECT 111.650 16.450 112.070 22.000 ;
        RECT 111.650 15.450 112.000 16.450 ;
        RECT 112.460 16.250 112.690 30.240 ;
        RECT 113.050 29.400 113.470 30.400 ;
        RECT 114.300 30.250 117.550 30.650 ;
        RECT 120.900 30.440 121.300 30.450 ;
        RECT 122.250 30.440 122.650 30.450 ;
        RECT 112.850 28.800 113.470 29.400 ;
        RECT 112.850 27.400 113.250 28.800 ;
        RECT 113.750 27.700 113.980 30.240 ;
        RECT 112.850 26.500 113.150 27.400 ;
        RECT 113.500 26.700 114.000 27.700 ;
        RECT 112.850 26.100 113.250 26.500 ;
        RECT 112.850 25.900 113.470 26.100 ;
        RECT 112.950 25.200 113.470 25.900 ;
        RECT 113.050 22.500 113.470 25.200 ;
        RECT 113.050 21.900 113.500 22.500 ;
        RECT 112.200 15.600 112.900 16.250 ;
        RECT 111.650 14.080 112.070 15.450 ;
        RECT 112.460 14.240 112.690 15.600 ;
        RECT 113.050 14.080 113.470 21.900 ;
        RECT 113.750 14.240 113.980 26.700 ;
        RECT 108.870 13.850 109.830 14.080 ;
        RECT 110.160 13.850 111.120 14.080 ;
        RECT 111.450 13.850 112.410 14.080 ;
        RECT 112.740 13.850 113.700 14.080 ;
        RECT 114.300 13.550 117.450 30.250 ;
        RECT 118.050 30.210 119.010 30.440 ;
        RECT 119.340 30.210 120.300 30.440 ;
        RECT 120.630 30.210 121.590 30.440 ;
        RECT 121.920 30.210 122.880 30.440 ;
        RECT 117.770 27.800 118.000 30.050 ;
        RECT 118.250 28.250 118.670 30.210 ;
        RECT 118.250 28.200 118.850 28.250 ;
        RECT 117.770 26.800 118.350 27.800 ;
        RECT 117.770 14.050 118.000 26.800 ;
        RECT 118.500 26.450 118.850 28.200 ;
        RECT 118.500 26.400 118.670 26.450 ;
        RECT 118.250 19.500 118.670 26.400 ;
        RECT 118.250 18.900 118.700 19.500 ;
        RECT 118.250 13.890 118.670 18.900 ;
        RECT 119.060 16.200 119.290 30.050 ;
        RECT 119.650 19.600 120.050 30.210 ;
        RECT 120.350 27.700 120.580 30.050 ;
        RECT 120.200 26.700 120.700 27.700 ;
        RECT 119.650 19.000 120.100 19.600 ;
        RECT 119.650 16.500 120.050 19.000 ;
        RECT 118.850 15.550 119.550 16.200 ;
        RECT 119.060 14.050 119.290 15.550 ;
        RECT 119.750 15.250 120.050 16.500 ;
        RECT 119.650 13.890 120.050 15.250 ;
        RECT 120.350 14.050 120.580 26.700 ;
        RECT 120.900 13.890 121.300 30.210 ;
        RECT 121.640 16.300 121.870 30.050 ;
        RECT 122.250 19.700 122.650 30.210 ;
        RECT 122.930 27.600 123.160 30.050 ;
        RECT 122.800 26.600 123.300 27.600 ;
        RECT 122.250 19.100 122.700 19.700 ;
        RECT 122.250 16.550 122.650 19.100 ;
        RECT 121.450 15.650 122.150 16.300 ;
        RECT 121.640 14.050 121.870 15.650 ;
        RECT 122.350 15.300 122.650 16.550 ;
        RECT 122.250 13.890 122.650 15.300 ;
        RECT 122.930 14.050 123.160 26.600 ;
        RECT 123.550 25.330 126.350 30.650 ;
        RECT 126.600 26.600 127.200 41.200 ;
        RECT 126.770 26.050 127.000 26.600 ;
        RECT 128.060 26.400 131.000 41.600 ;
        RECT 128.060 26.050 128.290 26.400 ;
        RECT 127.100 25.890 127.900 25.900 ;
        RECT 127.050 25.660 128.010 25.890 ;
        RECT 127.100 25.600 127.900 25.660 ;
        RECT 129.050 25.330 130.050 26.400 ;
        RECT 130.770 26.050 131.000 26.400 ;
        RECT 131.250 25.900 131.550 42.200 ;
        RECT 132.060 41.300 132.290 42.050 ;
        RECT 131.900 26.700 132.500 41.300 ;
        RECT 132.060 26.050 132.290 26.700 ;
        RECT 132.750 25.900 133.050 42.200 ;
        RECT 133.350 41.800 133.580 42.050 ;
        RECT 134.050 41.800 137.000 42.700 ;
        RECT 133.350 26.700 137.000 41.800 ;
        RECT 137.700 31.800 143.050 46.400 ;
        RECT 137.650 27.000 143.050 31.800 ;
        RECT 137.670 26.950 142.600 27.000 ;
        RECT 138.100 26.900 142.600 26.950 ;
        RECT 133.350 26.050 133.580 26.700 ;
        RECT 134.050 26.050 137.000 26.700 ;
        RECT 134.050 25.950 138.600 26.050 ;
        RECT 131.150 25.890 133.350 25.900 ;
        RECT 131.050 25.660 133.350 25.890 ;
        RECT 131.150 25.500 133.350 25.660 ;
        RECT 134.050 25.330 143.050 25.950 ;
        RECT 123.550 23.600 143.050 25.330 ;
        RECT 123.550 22.400 125.400 23.600 ;
        RECT 125.910 22.880 128.015 23.130 ;
        RECT 137.820 22.800 140.100 23.210 ;
        RECT 140.450 22.400 143.050 23.600 ;
        RECT 123.550 20.650 143.050 22.400 ;
        RECT 123.550 19.350 125.400 20.650 ;
        RECT 125.820 19.800 128.100 20.210 ;
        RECT 137.820 19.800 140.100 20.210 ;
        RECT 140.450 19.350 143.050 20.650 ;
        RECT 123.550 17.750 143.050 19.350 ;
        RECT 123.550 14.400 125.450 17.750 ;
        RECT 125.650 17.720 127.410 17.750 ;
        RECT 127.550 17.700 143.050 17.750 ;
        RECT 126.050 17.210 127.010 17.440 ;
        RECT 125.770 17.000 126.000 17.050 ;
        RECT 125.600 15.150 126.000 17.000 ;
        RECT 125.770 15.050 126.000 15.150 ;
        RECT 126.300 14.890 126.750 17.210 ;
        RECT 127.060 16.950 127.290 17.050 ;
        RECT 127.550 16.950 130.450 17.700 ;
        RECT 130.800 17.440 131.950 17.500 ;
        RECT 132.350 17.450 143.050 17.700 ;
        RECT 130.800 17.210 132.010 17.440 ;
        RECT 130.800 17.200 131.950 17.210 ;
        RECT 130.800 17.050 131.900 17.200 ;
        RECT 127.060 15.110 130.450 16.950 ;
        RECT 127.060 15.050 127.290 15.110 ;
        RECT 126.050 14.660 127.010 14.890 ;
        RECT 127.550 14.480 130.450 15.110 ;
        RECT 130.770 15.110 131.900 17.050 ;
        RECT 132.060 16.900 132.290 17.050 ;
        RECT 132.630 16.900 143.050 17.450 ;
        RECT 132.050 15.250 143.050 16.900 ;
        RECT 130.770 15.050 131.000 15.110 ;
        RECT 131.350 14.950 131.900 15.110 ;
        RECT 132.060 15.200 143.050 15.250 ;
        RECT 132.060 15.050 132.290 15.200 ;
        RECT 131.200 14.900 131.900 14.950 ;
        RECT 131.100 14.890 131.950 14.900 ;
        RECT 131.050 14.660 132.010 14.890 ;
        RECT 132.630 14.700 143.050 15.200 ;
        RECT 132.500 14.550 143.050 14.700 ;
        RECT 127.550 14.400 130.460 14.480 ;
        RECT 123.550 14.380 125.850 14.400 ;
        RECT 127.200 14.380 130.700 14.400 ;
        RECT 132.350 14.380 143.050 14.550 ;
        RECT 118.050 13.660 119.010 13.890 ;
        RECT 119.340 13.660 120.300 13.890 ;
        RECT 120.630 13.660 121.590 13.890 ;
        RECT 121.920 13.660 122.880 13.890 ;
        RECT 119.650 13.650 120.050 13.660 ;
        RECT 105.050 13.350 117.450 13.550 ;
        RECT 123.550 13.350 143.050 14.380 ;
        RECT 105.050 10.000 143.050 13.350 ;
      LAYER met2 ;
        RECT 98.600 207.650 99.500 208.300 ;
        RECT 97.950 206.450 98.550 207.100 ;
        RECT 121.950 205.840 122.450 210.070 ;
        RECT 123.550 208.450 124.050 210.070 ;
        RECT 123.500 207.490 124.050 208.450 ;
        RECT 123.465 207.210 124.050 207.490 ;
        RECT 123.500 207.200 124.050 207.210 ;
        RECT 82.970 204.850 83.730 205.550 ;
        RECT 83.000 141.075 86.000 204.850 ;
        RECT 94.300 203.900 95.300 205.100 ;
        RECT 96.025 204.660 97.085 205.660 ;
        RECT 110.050 205.340 122.450 205.840 ;
        RECT 96.055 203.500 97.055 204.660 ;
        RECT 96.010 202.500 97.100 203.500 ;
        RECT 91.205 201.610 91.505 201.640 ;
        RECT 94.405 201.610 100.055 201.860 ;
        RECT 91.205 201.310 100.055 201.610 ;
        RECT 91.205 201.280 91.505 201.310 ;
        RECT 99.605 201.210 100.005 201.310 ;
        RECT 92.905 199.160 97.355 201.010 ;
        RECT 90.255 196.260 96.555 197.660 ;
        RECT 91.755 195.360 92.155 195.410 ;
        RECT 94.555 195.360 94.955 195.410 ;
        RECT 91.755 195.060 94.955 195.360 ;
        RECT 91.755 195.010 92.155 195.060 ;
        RECT 94.555 195.010 94.955 195.060 ;
        RECT 94.555 190.460 94.955 190.660 ;
        RECT 94.505 189.860 94.955 190.460 ;
        RECT 94.555 189.760 94.955 189.860 ;
        RECT 98.055 189.760 98.555 189.860 ;
        RECT 94.555 189.460 98.555 189.760 ;
        RECT 91.755 185.110 92.155 185.160 ;
        RECT 94.405 185.110 94.955 185.160 ;
        RECT 91.755 184.810 95.005 185.110 ;
        RECT 91.755 184.760 92.155 184.810 ;
        RECT 94.605 184.760 94.955 184.810 ;
        RECT 90.955 184.560 91.255 184.590 ;
        RECT 90.955 184.260 91.405 184.560 ;
        RECT 95.405 184.260 95.855 184.560 ;
        RECT 90.955 183.760 91.355 184.260 ;
        RECT 95.455 183.760 95.855 184.260 ;
        RECT 99.555 183.760 100.105 183.910 ;
        RECT 90.955 183.410 100.105 183.760 ;
        RECT 99.555 183.260 100.105 183.410 ;
        RECT 110.050 162.690 110.550 205.340 ;
        RECT 123.550 204.840 124.050 207.200 ;
        RECT 111.050 204.340 124.050 204.840 ;
        RECT 111.050 174.690 111.550 204.340 ;
        RECT 124.450 203.640 124.950 210.070 ;
        RECT 112.050 203.140 124.950 203.640 ;
        RECT 112.050 186.690 112.550 203.140 ;
        RECT 125.450 202.840 125.950 210.070 ;
        RECT 113.150 202.340 125.950 202.840 ;
        RECT 126.650 202.940 127.150 215.850 ;
        RECT 127.650 203.940 128.150 218.150 ;
        RECT 128.650 205.140 129.150 215.800 ;
        RECT 129.750 205.940 130.250 215.750 ;
        RECT 131.800 205.940 135.200 205.950 ;
        RECT 129.750 205.440 142.500 205.940 ;
        RECT 131.800 205.140 135.200 205.150 ;
        RECT 128.650 204.640 141.550 205.140 ;
        RECT 131.800 204.630 135.200 204.640 ;
        RECT 127.650 203.440 140.650 203.940 ;
        RECT 126.650 202.440 139.550 202.940 ;
        RECT 113.150 198.790 113.650 202.340 ;
        RECT 115.195 201.990 135.905 201.995 ;
        RECT 115.195 201.590 136.800 201.990 ;
        RECT 138.550 201.640 139.550 202.440 ;
        RECT 115.195 201.585 135.905 201.590 ;
        RECT 115.300 201.190 116.100 201.585 ;
        RECT 136.170 201.190 136.800 201.590 ;
        RECT 115.200 200.190 116.200 201.190 ;
        RECT 113.000 198.090 113.700 198.790 ;
        RECT 115.500 195.090 116.000 200.190 ;
        RECT 118.200 199.290 119.500 201.190 ;
        RECT 117.800 198.990 119.500 199.290 ;
        RECT 120.100 199.840 123.400 200.290 ;
        RECT 117.800 198.940 119.100 198.990 ;
        RECT 117.050 198.090 117.450 198.790 ;
        RECT 120.100 197.990 120.600 199.840 ;
        RECT 117.700 197.390 120.600 197.990 ;
        RECT 120.850 196.990 122.650 197.590 ;
        RECT 120.850 195.090 121.350 196.990 ;
        RECT 122.800 196.790 123.200 199.690 ;
        RECT 122.000 196.190 124.100 196.790 ;
        RECT 115.500 194.490 121.350 195.090 ;
        RECT 115.500 194.390 116.000 194.490 ;
        RECT 122.800 193.990 123.200 196.190 ;
        RECT 122.100 193.390 124.100 193.990 ;
        RECT 115.500 190.190 116.000 191.990 ;
        RECT 116.500 191.090 122.100 191.590 ;
        RECT 122.800 191.090 123.200 193.390 ;
        RECT 116.500 190.490 124.000 191.090 ;
        RECT 116.500 190.390 122.100 190.490 ;
        RECT 120.700 190.190 122.100 190.390 ;
        RECT 115.200 188.190 116.200 190.190 ;
        RECT 113.000 186.690 113.600 186.790 ;
        RECT 112.050 186.190 113.600 186.690 ;
        RECT 113.000 186.090 113.600 186.190 ;
        RECT 115.500 183.090 116.000 188.190 ;
        RECT 118.200 187.290 119.500 189.190 ;
        RECT 117.800 186.990 119.500 187.290 ;
        RECT 120.100 187.840 123.400 188.290 ;
        RECT 117.800 186.940 119.100 186.990 ;
        RECT 117.050 186.090 117.450 186.790 ;
        RECT 120.100 185.990 120.600 187.840 ;
        RECT 117.700 185.390 120.600 185.990 ;
        RECT 120.850 184.990 122.650 185.590 ;
        RECT 120.850 183.090 121.350 184.990 ;
        RECT 122.800 184.790 123.200 187.690 ;
        RECT 122.000 184.190 124.100 184.790 ;
        RECT 115.500 182.490 121.350 183.090 ;
        RECT 115.500 182.390 116.000 182.490 ;
        RECT 122.800 181.990 123.200 184.190 ;
        RECT 122.100 181.390 124.100 181.990 ;
        RECT 115.500 178.190 116.000 179.990 ;
        RECT 116.500 179.090 122.100 179.590 ;
        RECT 122.800 179.090 123.200 181.390 ;
        RECT 116.500 178.490 124.000 179.090 ;
        RECT 116.500 178.390 122.100 178.490 ;
        RECT 120.700 178.190 122.100 178.390 ;
        RECT 115.200 176.190 116.200 178.190 ;
        RECT 113.075 174.690 113.525 174.710 ;
        RECT 111.050 174.190 113.550 174.690 ;
        RECT 113.075 174.170 113.525 174.190 ;
        RECT 115.500 171.090 116.000 176.190 ;
        RECT 118.200 175.290 119.500 177.190 ;
        RECT 117.800 174.990 119.500 175.290 ;
        RECT 120.100 175.840 123.400 176.290 ;
        RECT 117.800 174.940 119.100 174.990 ;
        RECT 117.050 174.090 117.450 174.790 ;
        RECT 120.100 173.990 120.600 175.840 ;
        RECT 117.700 173.390 120.600 173.990 ;
        RECT 120.850 172.990 122.650 173.590 ;
        RECT 120.850 171.090 121.350 172.990 ;
        RECT 122.800 172.790 123.200 175.690 ;
        RECT 122.000 172.190 124.100 172.790 ;
        RECT 115.500 170.490 121.350 171.090 ;
        RECT 115.500 170.390 116.000 170.490 ;
        RECT 122.800 169.990 123.200 172.190 ;
        RECT 122.100 169.390 124.100 169.990 ;
        RECT 115.500 166.190 116.000 167.990 ;
        RECT 116.500 167.090 122.100 167.590 ;
        RECT 122.800 167.090 123.200 169.390 ;
        RECT 116.500 166.490 124.000 167.090 ;
        RECT 116.500 166.390 122.100 166.490 ;
        RECT 120.700 166.190 122.100 166.390 ;
        RECT 115.200 164.190 116.200 166.190 ;
        RECT 113.175 162.690 113.625 162.710 ;
        RECT 110.050 162.190 113.650 162.690 ;
        RECT 113.175 162.170 113.625 162.190 ;
        RECT 115.500 159.090 116.000 164.190 ;
        RECT 118.200 163.290 119.500 165.190 ;
        RECT 117.800 162.990 119.500 163.290 ;
        RECT 120.100 163.840 123.400 164.290 ;
        RECT 117.800 162.940 119.100 162.990 ;
        RECT 117.050 162.090 117.450 162.790 ;
        RECT 120.100 161.990 120.600 163.840 ;
        RECT 117.700 161.390 120.600 161.990 ;
        RECT 120.850 160.990 122.650 161.590 ;
        RECT 120.850 159.090 121.350 160.990 ;
        RECT 122.800 160.790 123.200 163.690 ;
        RECT 122.000 160.190 124.100 160.790 ;
        RECT 115.500 158.490 121.350 159.090 ;
        RECT 115.500 158.390 116.000 158.490 ;
        RECT 122.800 157.990 123.200 160.190 ;
        RECT 122.100 157.390 124.100 157.990 ;
        RECT 115.500 154.190 116.000 155.990 ;
        RECT 116.500 155.090 122.100 155.590 ;
        RECT 122.800 155.090 123.200 157.390 ;
        RECT 116.500 154.490 124.000 155.090 ;
        RECT 116.500 154.390 122.100 154.490 ;
        RECT 120.700 154.190 122.100 154.390 ;
        RECT 115.000 152.690 116.500 154.190 ;
        RECT 110.500 150.450 111.500 151.550 ;
        RECT 112.000 149.000 113.000 149.550 ;
        RECT 115.240 149.000 116.410 152.690 ;
        RECT 125.000 151.690 127.000 201.190 ;
        RECT 135.800 200.190 136.800 201.190 ;
        RECT 129.900 199.990 131.300 200.190 ;
        RECT 129.900 199.890 135.500 199.990 ;
        RECT 128.000 199.290 135.500 199.890 ;
        RECT 128.800 196.990 129.200 199.290 ;
        RECT 129.900 198.790 135.500 199.290 ;
        RECT 136.000 198.390 136.500 200.190 ;
        RECT 127.900 196.390 129.900 196.990 ;
        RECT 128.800 194.190 129.200 196.390 ;
        RECT 136.000 195.890 136.500 195.990 ;
        RECT 130.650 195.290 136.500 195.890 ;
        RECT 127.900 193.590 130.000 194.190 ;
        RECT 128.800 190.690 129.200 193.590 ;
        RECT 130.650 193.390 131.150 195.290 ;
        RECT 129.350 192.790 131.150 193.390 ;
        RECT 131.400 192.390 134.300 192.990 ;
        RECT 131.400 190.540 131.900 192.390 ;
        RECT 134.550 191.590 134.950 192.290 ;
        RECT 132.900 191.390 134.200 191.440 ;
        RECT 128.600 190.090 131.900 190.540 ;
        RECT 132.500 191.090 134.200 191.390 ;
        RECT 132.500 189.190 133.800 191.090 ;
        RECT 136.000 190.190 136.500 195.290 ;
        RECT 139.050 192.290 139.550 201.640 ;
        RECT 138.500 191.490 139.600 192.290 ;
        RECT 135.800 188.190 136.800 190.190 ;
        RECT 129.900 187.990 131.300 188.190 ;
        RECT 129.900 187.890 135.500 187.990 ;
        RECT 128.000 187.290 135.500 187.890 ;
        RECT 128.800 184.990 129.200 187.290 ;
        RECT 129.900 186.790 135.500 187.290 ;
        RECT 136.000 186.390 136.500 188.190 ;
        RECT 127.900 184.390 129.900 184.990 ;
        RECT 128.800 182.190 129.200 184.390 ;
        RECT 136.000 183.890 136.500 183.990 ;
        RECT 130.650 183.290 136.500 183.890 ;
        RECT 127.900 181.590 130.000 182.190 ;
        RECT 128.800 178.690 129.200 181.590 ;
        RECT 130.650 181.390 131.150 183.290 ;
        RECT 129.350 180.790 131.150 181.390 ;
        RECT 131.400 180.390 134.300 180.990 ;
        RECT 131.400 178.540 131.900 180.390 ;
        RECT 134.550 179.590 134.950 180.290 ;
        RECT 132.900 179.390 134.200 179.440 ;
        RECT 128.600 178.090 131.900 178.540 ;
        RECT 132.500 179.090 134.200 179.390 ;
        RECT 132.500 177.190 133.800 179.090 ;
        RECT 136.000 178.190 136.500 183.290 ;
        RECT 140.150 180.140 140.650 203.440 ;
        RECT 138.550 179.640 140.650 180.140 ;
        RECT 135.800 176.190 136.800 178.190 ;
        RECT 129.900 175.990 131.300 176.190 ;
        RECT 129.900 175.890 135.500 175.990 ;
        RECT 128.000 175.290 135.500 175.890 ;
        RECT 128.800 172.990 129.200 175.290 ;
        RECT 129.900 174.790 135.500 175.290 ;
        RECT 136.000 174.390 136.500 176.190 ;
        RECT 127.900 172.390 129.900 172.990 ;
        RECT 128.800 170.190 129.200 172.390 ;
        RECT 136.000 171.890 136.500 171.990 ;
        RECT 130.650 171.290 136.500 171.890 ;
        RECT 127.900 169.590 130.000 170.190 ;
        RECT 128.800 166.690 129.200 169.590 ;
        RECT 130.650 169.390 131.150 171.290 ;
        RECT 129.350 168.790 131.150 169.390 ;
        RECT 131.400 168.390 134.300 168.990 ;
        RECT 131.400 166.540 131.900 168.390 ;
        RECT 134.550 167.590 134.950 168.290 ;
        RECT 132.900 167.390 134.200 167.440 ;
        RECT 128.600 166.090 131.900 166.540 ;
        RECT 132.500 167.090 134.200 167.390 ;
        RECT 132.500 165.190 133.800 167.090 ;
        RECT 136.000 166.190 136.500 171.290 ;
        RECT 141.050 168.140 141.550 204.640 ;
        RECT 138.505 167.640 141.550 168.140 ;
        RECT 141.050 167.590 141.550 167.640 ;
        RECT 135.800 164.190 136.800 166.190 ;
        RECT 129.900 163.990 131.300 164.190 ;
        RECT 129.900 163.890 135.500 163.990 ;
        RECT 128.000 163.290 135.500 163.890 ;
        RECT 128.800 160.990 129.200 163.290 ;
        RECT 129.900 162.790 135.500 163.290 ;
        RECT 136.000 162.390 136.500 164.190 ;
        RECT 127.900 160.390 129.900 160.990 ;
        RECT 128.800 158.190 129.200 160.390 ;
        RECT 136.000 159.890 136.500 159.990 ;
        RECT 130.650 159.290 136.500 159.890 ;
        RECT 127.900 157.590 130.000 158.190 ;
        RECT 128.800 154.690 129.200 157.590 ;
        RECT 130.650 157.390 131.150 159.290 ;
        RECT 129.350 156.790 131.150 157.390 ;
        RECT 131.400 156.390 134.300 156.990 ;
        RECT 131.400 154.540 131.900 156.390 ;
        RECT 134.550 155.590 134.950 156.290 ;
        RECT 132.900 155.390 134.200 155.440 ;
        RECT 128.600 154.090 131.900 154.540 ;
        RECT 132.500 155.090 134.200 155.390 ;
        RECT 132.500 153.190 133.800 155.090 ;
        RECT 136.000 154.190 136.500 159.290 ;
        RECT 138.505 155.990 140.600 156.140 ;
        RECT 142.050 156.015 142.500 205.440 ;
        RECT 141.800 155.990 142.500 156.015 ;
        RECT 138.505 155.640 142.500 155.990 ;
        RECT 138.575 155.590 142.500 155.640 ;
        RECT 138.575 155.565 141.000 155.590 ;
        RECT 135.500 152.690 137.000 154.190 ;
        RECT 125.400 150.390 126.200 151.690 ;
        RECT 126.900 150.490 129.900 150.590 ;
        RECT 125.300 149.090 126.400 150.390 ;
        RECT 126.750 150.090 130.550 150.490 ;
        RECT 111.000 148.450 113.000 149.000 ;
        RECT 111.000 147.550 112.000 148.450 ;
        RECT 110.500 146.450 112.000 147.550 ;
        RECT 82.980 138.125 86.020 141.075 ;
        RECT 83.000 138.100 86.000 138.125 ;
        RECT 111.000 133.000 112.000 146.450 ;
        RECT 115.000 145.000 117.000 149.000 ;
        RECT 115.000 133.475 116.000 145.000 ;
        RECT 126.900 138.055 129.900 150.090 ;
        RECT 133.000 150.000 135.000 152.500 ;
        RECT 135.700 148.490 136.900 152.690 ;
        RECT 135.600 146.190 136.900 148.490 ;
        RECT 136.070 145.000 136.670 146.190 ;
        RECT 111.150 128.820 111.950 133.000 ;
        RECT 113.300 132.925 116.025 133.475 ;
        RECT 113.300 119.800 113.850 132.925 ;
        RECT 106.500 62.950 108.000 64.550 ;
        RECT 111.000 62.950 112.500 64.550 ;
        RECT 119.950 61.000 120.450 61.050 ;
        RECT 122.650 61.000 123.650 62.200 ;
        RECT 125.950 61.000 126.450 61.050 ;
        RECT 128.750 61.000 129.750 62.400 ;
        RECT 131.950 61.000 132.450 61.050 ;
        RECT 119.550 60.000 123.650 61.000 ;
        RECT 125.550 60.000 133.050 61.000 ;
        RECT 119.950 59.950 120.450 60.000 ;
        RECT 119.950 58.500 120.450 58.550 ;
        RECT 122.650 58.500 123.650 60.000 ;
        RECT 125.950 59.950 126.450 60.000 ;
        RECT 125.950 58.500 126.450 58.550 ;
        RECT 128.750 58.500 129.750 60.000 ;
        RECT 131.950 59.950 132.450 60.000 ;
        RECT 131.950 58.500 132.450 58.550 ;
        RECT 119.550 57.500 123.650 58.500 ;
        RECT 125.550 57.500 133.050 58.500 ;
        RECT 119.950 57.450 120.450 57.500 ;
        RECT 119.950 56.500 120.450 56.550 ;
        RECT 122.650 56.500 123.650 57.500 ;
        RECT 125.950 57.450 126.450 57.500 ;
        RECT 128.750 56.500 129.750 57.500 ;
        RECT 131.950 57.450 132.450 57.500 ;
        RECT 131.950 56.500 132.450 56.550 ;
        RECT 119.550 55.500 123.650 56.500 ;
        RECT 125.550 55.500 133.050 56.500 ;
        RECT 119.950 55.450 120.450 55.500 ;
        RECT 119.950 54.000 120.450 54.050 ;
        RECT 122.650 54.000 123.650 55.500 ;
        RECT 125.950 54.000 126.450 54.050 ;
        RECT 128.750 54.000 129.750 55.500 ;
        RECT 131.950 55.450 132.450 55.500 ;
        RECT 131.950 54.000 132.450 54.050 ;
        RECT 119.550 53.000 123.650 54.000 ;
        RECT 125.550 53.000 133.050 54.000 ;
        RECT 119.950 52.950 120.450 53.000 ;
        RECT 122.650 50.750 123.650 53.000 ;
        RECT 125.950 52.950 126.450 53.000 ;
        RECT 128.750 50.750 129.750 53.000 ;
        RECT 131.950 52.950 132.450 53.000 ;
        RECT 106.550 50.500 107.550 50.550 ;
        RECT 125.350 50.500 125.750 50.550 ;
        RECT 126.550 50.500 126.950 50.550 ;
        RECT 131.350 50.500 131.750 50.550 ;
        RECT 132.550 50.500 132.950 50.550 ;
        RECT 105.050 49.500 135.050 50.500 ;
        RECT 106.550 49.450 107.550 49.500 ;
        RECT 114.950 49.450 115.350 49.500 ;
        RECT 125.350 49.450 125.750 49.500 ;
        RECT 126.550 49.450 126.950 49.500 ;
        RECT 131.350 49.450 131.750 49.500 ;
        RECT 132.550 49.450 132.950 49.500 ;
        RECT 105.050 48.500 106.050 48.550 ;
        RECT 109.250 48.500 109.550 48.550 ;
        RECT 119.250 48.500 119.750 48.550 ;
        RECT 120.550 48.500 121.050 48.550 ;
        RECT 105.050 47.500 135.050 48.500 ;
        RECT 105.050 47.450 106.050 47.500 ;
        RECT 109.250 47.450 109.550 47.500 ;
        RECT 119.250 47.450 119.750 47.500 ;
        RECT 120.550 47.450 121.050 47.500 ;
        RECT 137.550 44.900 143.050 45.500 ;
        RECT 122.650 44.800 123.650 44.850 ;
        RECT 124.650 44.800 125.650 44.850 ;
        RECT 126.450 44.800 127.450 44.850 ;
        RECT 122.650 43.800 127.450 44.800 ;
        RECT 122.650 43.750 123.650 43.800 ;
        RECT 124.650 43.750 125.650 43.800 ;
        RECT 106.550 42.000 107.550 42.050 ;
        RECT 105.050 41.000 125.550 42.000 ;
        RECT 106.550 40.950 107.550 41.000 ;
        RECT 123.050 40.950 123.350 41.000 ;
        RECT 105.050 40.500 106.050 40.550 ;
        RECT 117.750 40.500 118.050 40.550 ;
        RECT 105.050 39.500 125.550 40.500 ;
        RECT 105.050 39.450 106.050 39.500 ;
        RECT 117.750 39.450 118.050 39.500 ;
        RECT 102.155 38.000 125.550 39.000 ;
        RECT 99.950 36.500 125.550 37.500 ;
        RECT 107.050 35.000 115.550 36.000 ;
        RECT 116.550 35.000 125.550 36.000 ;
        RECT 110.550 28.500 112.050 35.000 ;
        RECT 119.550 28.500 121.050 35.000 ;
        RECT 107.550 26.500 115.550 28.500 ;
        RECT 116.550 26.500 124.550 28.500 ;
        RECT 126.450 26.600 127.450 43.800 ;
        RECT 128.650 43.400 143.050 44.900 ;
        RECT 131.750 26.800 132.750 43.400 ;
        RECT 137.550 43.000 143.050 43.400 ;
        RECT 137.750 29.580 143.150 30.800 ;
        RECT 126.950 25.400 133.650 26.200 ;
        RECT 125.650 23.550 128.200 24.050 ;
        RECT 98.250 21.500 123.050 23.000 ;
        RECT 98.250 5.000 99.750 21.500 ;
        RECT 101.200 18.500 123.050 20.000 ;
        RECT 125.600 18.850 128.200 23.550 ;
        RECT 101.200 6.105 102.700 18.500 ;
        RECT 125.600 18.350 128.150 18.850 ;
        RECT 137.700 18.800 143.150 29.580 ;
        RECT 137.700 18.750 140.300 18.800 ;
        RECT 126.050 17.550 127.550 18.350 ;
        RECT 125.650 17.000 125.950 17.050 ;
        RECT 107.050 16.450 123.550 17.000 ;
        RECT 124.550 16.450 126.000 17.000 ;
        RECT 107.050 15.350 126.000 16.450 ;
        RECT 107.050 15.000 123.550 15.350 ;
        RECT 124.550 15.150 126.000 15.350 ;
        RECT 126.300 16.500 127.550 17.550 ;
        RECT 125.650 15.100 125.950 15.150 ;
        RECT 126.300 15.000 131.800 16.500 ;
        RECT 126.300 14.500 127.550 15.000 ;
        RECT 109.000 10.950 113.000 12.050 ;
        RECT 121.500 10.450 124.500 12.050 ;
        RECT 97.650 3.100 100.000 5.000 ;
      LAYER met3 ;
        RECT 46.655 220.760 48.145 220.785 ;
        RECT 3.550 219.260 48.150 220.760 ;
        RECT 51.855 220.750 53.345 220.775 ;
        RECT 51.850 220.730 82.150 220.750 ;
        RECT 82.450 220.730 83.450 220.750 ;
        RECT 46.655 219.235 48.145 219.260 ;
        RECT 51.850 219.250 83.450 220.730 ;
        RECT 100.650 219.495 116.050 219.500 ;
        RECT 51.855 219.225 53.345 219.250 ;
        RECT 81.600 219.160 82.600 219.250 ;
        RECT 100.625 218.505 116.050 219.495 ;
        RECT 100.650 218.500 116.050 218.505 ;
        RECT 127.550 217.500 128.250 218.350 ;
        RECT 102.205 216.700 103.195 216.725 ;
        RECT 102.200 215.700 119.250 216.700 ;
        RECT 102.205 215.675 103.195 215.700 ;
        RECT 121.740 213.200 122.060 213.240 ;
        RECT 129.885 213.200 130.215 213.215 ;
        RECT 121.740 212.900 130.215 213.200 ;
        RECT 121.740 212.860 122.060 212.900 ;
        RECT 129.885 212.885 130.215 212.900 ;
        RECT 125.390 211.500 125.770 211.510 ;
        RECT 128.785 211.500 129.115 211.515 ;
        RECT 125.390 211.200 129.115 211.500 ;
        RECT 125.390 211.190 125.770 211.200 ;
        RECT 128.785 211.185 129.115 211.200 ;
        RECT 126.685 210.100 127.015 210.115 ;
        RECT 132.780 210.100 133.100 210.140 ;
        RECT 126.685 209.800 133.100 210.100 ;
        RECT 126.685 209.785 127.015 209.800 ;
        RECT 132.780 209.760 133.100 209.800 ;
        RECT 125.485 209.200 125.815 209.215 ;
        RECT 136.460 209.200 136.780 209.240 ;
        RECT 125.485 208.900 136.780 209.200 ;
        RECT 125.485 208.885 125.815 208.900 ;
        RECT 136.460 208.860 136.780 208.900 ;
        RECT 124.485 208.300 124.815 208.315 ;
        RECT 140.140 208.300 140.460 208.340 ;
        RECT 98.600 208.150 99.500 208.300 ;
        RECT 88.420 207.750 99.500 208.150 ;
        RECT 124.485 208.000 140.460 208.300 ;
        RECT 124.485 207.985 124.815 208.000 ;
        RECT 140.140 207.960 140.460 208.000 ;
        RECT 98.600 207.650 99.500 207.750 ;
        RECT 123.485 207.500 123.815 207.515 ;
        RECT 143.790 207.500 144.170 207.510 ;
        RECT 123.485 207.200 144.170 207.500 ;
        RECT 123.485 207.185 123.815 207.200 ;
        RECT 143.790 207.190 144.170 207.200 ;
        RECT 98.030 206.900 98.480 206.925 ;
        RECT 84.850 206.500 98.480 206.900 ;
        RECT 121.935 206.850 122.265 206.865 ;
        RECT 147.500 206.850 147.820 206.890 ;
        RECT 121.935 206.550 147.820 206.850 ;
        RECT 121.935 206.535 122.265 206.550 ;
        RECT 147.500 206.510 147.820 206.550 ;
        RECT 98.030 206.475 98.480 206.500 ;
        RECT 4.100 204.750 7.600 205.500 ;
        RECT 94.430 204.750 95.180 204.775 ;
        RECT 4.100 204.050 95.180 204.750 ;
        RECT 4.100 202.300 7.600 204.050 ;
        RECT 94.430 204.025 95.180 204.050 ;
        RECT 96.030 203.500 97.080 203.525 ;
        RECT 53.970 202.500 97.080 203.500 ;
        RECT 96.030 202.475 97.080 202.500 ;
        RECT 118.000 199.690 127.000 201.190 ;
        RECT 125.000 199.190 127.000 199.690 ;
        RECT 113.000 198.690 113.500 198.790 ;
        RECT 116.500 198.690 117.500 199.190 ;
        RECT 113.000 198.190 117.500 198.690 ;
        RECT 113.000 198.090 113.500 198.190 ;
        RECT 116.500 197.690 117.500 198.190 ;
        RECT 134.500 192.190 135.500 192.690 ;
        RECT 138.500 192.190 139.000 192.290 ;
        RECT 134.500 192.140 139.000 192.190 ;
        RECT 134.500 191.690 139.025 192.140 ;
        RECT 134.500 191.190 135.500 191.690 ;
        RECT 138.500 191.640 139.025 191.690 ;
        RECT 138.500 191.590 139.000 191.640 ;
        RECT 125.000 189.190 134.000 190.690 ;
        RECT 118.000 187.690 127.000 189.190 ;
        RECT 113.000 186.690 113.500 186.790 ;
        RECT 116.500 186.690 117.500 187.190 ;
        RECT 113.000 186.190 117.500 186.690 ;
        RECT 113.000 186.090 113.500 186.190 ;
        RECT 116.500 185.690 117.500 186.190 ;
        RECT 134.500 180.190 135.500 180.690 ;
        RECT 138.500 180.190 139.000 180.290 ;
        RECT 134.500 180.140 139.000 180.190 ;
        RECT 134.500 179.690 139.025 180.140 ;
        RECT 134.500 179.190 135.500 179.690 ;
        RECT 138.500 179.640 139.025 179.690 ;
        RECT 138.500 179.590 139.000 179.640 ;
        RECT 125.000 177.190 134.000 178.690 ;
        RECT 118.000 175.690 127.000 177.190 ;
        RECT 113.000 174.690 113.500 174.790 ;
        RECT 116.500 174.690 117.500 175.190 ;
        RECT 113.000 174.190 117.500 174.690 ;
        RECT 113.000 174.090 113.500 174.190 ;
        RECT 116.500 173.690 117.500 174.190 ;
        RECT 134.500 168.190 135.500 168.690 ;
        RECT 138.500 168.190 139.000 168.290 ;
        RECT 134.500 168.165 139.000 168.190 ;
        RECT 134.500 167.690 139.075 168.165 ;
        RECT 134.500 167.190 135.500 167.690 ;
        RECT 138.500 167.615 139.075 167.690 ;
        RECT 138.500 167.590 139.000 167.615 ;
        RECT 125.000 165.190 134.000 166.690 ;
        RECT 118.000 163.690 127.000 165.190 ;
        RECT 113.000 162.690 113.500 162.790 ;
        RECT 116.500 162.690 117.500 163.190 ;
        RECT 113.000 162.190 117.500 162.690 ;
        RECT 113.000 162.090 113.500 162.190 ;
        RECT 116.500 161.690 117.500 162.190 ;
        RECT 52.755 160.250 54.245 160.275 ;
        RECT 52.500 158.750 107.280 160.250 ;
        RECT 52.755 158.725 54.245 158.750 ;
        RECT 134.500 156.190 135.500 156.690 ;
        RECT 138.500 156.190 139.000 156.290 ;
        RECT 134.500 156.165 139.000 156.190 ;
        RECT 134.500 155.690 139.075 156.165 ;
        RECT 134.500 155.190 135.500 155.690 ;
        RECT 138.500 155.615 139.075 155.690 ;
        RECT 138.500 155.590 139.000 155.615 ;
        RECT 125.000 154.690 127.000 155.190 ;
        RECT 125.000 153.190 134.000 154.690 ;
        RECT 4.755 147.750 6.245 147.775 ;
        RECT 110.000 147.750 114.000 152.000 ;
        RECT 133.000 150.000 135.000 152.500 ;
        RECT 4.750 146.250 114.000 147.750 ;
        RECT 4.755 146.225 6.245 146.250 ;
        RECT 110.000 146.000 114.000 146.250 ;
        RECT 126.875 141.100 129.925 141.125 ;
        RECT 83.000 138.100 129.925 141.100 ;
        RECT 126.875 138.075 129.925 138.100 ;
        RECT 89.700 120.000 114.200 121.000 ;
        RECT 4.255 64.250 5.745 64.275 ;
        RECT 105.500 64.250 115.500 66.500 ;
        RECT 4.250 62.750 115.500 64.250 ;
        RECT 4.255 62.725 5.745 62.750 ;
        RECT 105.500 61.000 115.500 62.750 ;
        RECT 141.250 44.500 157.150 44.850 ;
        RECT 141.250 44.495 157.160 44.500 ;
        RECT 141.250 43.905 157.185 44.495 ;
        RECT 141.250 43.900 157.160 43.905 ;
        RECT 141.250 43.850 157.150 43.900 ;
        RECT 141.250 43.800 155.800 43.850 ;
        RECT 102.050 37.900 103.350 39.100 ;
        RECT 100.550 36.400 101.750 37.650 ;
        RECT 105.050 12.450 127.000 12.500 ;
        RECT 52.705 12.100 54.195 12.125 ;
        RECT 105.050 12.100 127.300 12.450 ;
        RECT 52.700 10.600 127.300 12.100 ;
        RECT 52.705 10.575 54.195 10.600 ;
        RECT 105.050 10.000 127.300 10.600 ;
        RECT 119.500 9.750 127.300 10.000 ;
        RECT 101.175 7.650 102.725 7.675 ;
        RECT 101.175 6.150 136.700 7.650 ;
        RECT 101.175 6.125 102.725 6.150 ;
        RECT 98.225 4.850 99.775 4.875 ;
        RECT 98.225 3.350 114.050 4.850 ;
        RECT 98.225 3.325 99.775 3.350 ;
      LAYER met4 ;
        RECT 33.730 224.760 37.110 225.060 ;
        RECT 37.410 224.760 40.790 225.060 ;
        RECT 41.090 224.760 44.470 225.060 ;
        RECT 44.770 224.760 48.150 225.060 ;
        RECT 48.450 224.760 51.830 225.060 ;
        RECT 52.130 224.760 55.510 225.060 ;
        RECT 55.810 224.760 59.190 225.060 ;
        RECT 3.990 220.065 4.290 224.760 ;
        RECT 7.670 220.065 7.970 224.760 ;
        RECT 11.350 220.165 11.650 224.760 ;
        RECT 15.030 220.165 15.330 224.760 ;
        RECT 3.975 219.735 4.305 220.065 ;
        RECT 7.655 219.735 7.985 220.065 ;
        RECT 11.335 219.835 11.665 220.165 ;
        RECT 15.015 219.835 15.345 220.165 ;
        RECT 18.710 220.065 19.010 224.760 ;
        RECT 22.390 220.165 22.690 224.760 ;
        RECT 26.070 220.165 26.370 224.760 ;
        RECT 29.750 220.165 30.050 224.760 ;
        RECT 18.695 219.735 19.025 220.065 ;
        RECT 22.375 219.835 22.705 220.165 ;
        RECT 26.055 219.835 26.385 220.165 ;
        RECT 29.735 219.835 30.065 220.165 ;
        RECT 33.450 220.065 33.750 224.760 ;
        RECT 33.435 219.735 33.765 220.065 ;
        RECT 46.650 219.260 49.000 220.760 ;
        RECT 50.500 219.250 53.350 220.750 ;
        RECT 62.870 220.165 63.170 224.760 ;
        RECT 66.550 220.165 66.850 224.760 ;
        RECT 70.230 220.165 70.530 224.760 ;
        RECT 73.910 220.165 74.210 224.760 ;
        RECT 77.590 220.165 77.890 224.760 ;
        RECT 62.855 219.835 63.185 220.165 ;
        RECT 66.535 219.835 66.865 220.165 ;
        RECT 70.215 219.835 70.545 220.165 ;
        RECT 73.895 219.835 74.225 220.165 ;
        RECT 77.575 219.835 77.905 220.165 ;
        RECT 81.270 220.065 81.570 224.760 ;
        RECT 81.255 219.735 81.585 220.065 ;
        RECT 84.950 206.865 85.250 224.760 ;
        RECT 88.630 212.400 88.930 224.760 ;
        RECT 88.450 211.700 89.150 212.400 ;
        RECT 88.450 208.155 88.850 211.700 ;
        RECT 88.445 207.745 88.855 208.155 ;
        RECT 84.935 206.535 85.265 206.865 ;
        RECT 4.100 204.850 7.600 205.500 ;
        RECT 2.500 203.350 7.600 204.850 ;
        RECT 53.995 203.500 55.005 203.505 ;
        RECT 4.100 202.300 7.600 203.350 ;
        RECT 50.500 202.500 55.005 203.500 ;
        RECT 53.995 202.495 55.005 202.500 ;
        RECT 50.500 158.750 54.250 160.250 ;
        RECT 2.500 146.250 6.250 147.750 ;
        RECT 89.895 119.995 90.905 121.005 ;
        RECT 2.500 62.750 5.750 64.250 ;
        RECT 50.500 10.600 54.200 12.100 ;
        RECT 89.900 3.500 90.900 119.995 ;
        RECT 100.650 37.530 101.650 219.500 ;
        RECT 114.390 219.115 114.690 224.760 ;
        RECT 114.375 218.785 114.705 219.115 ;
        RECT 102.200 39.030 103.200 216.700 ;
        RECT 118.070 216.165 118.370 224.760 ;
        RECT 118.055 215.835 118.385 216.165 ;
        RECT 121.750 213.215 122.050 224.760 ;
        RECT 121.735 212.885 122.065 213.215 ;
        RECT 125.430 211.515 125.730 224.760 ;
        RECT 127.785 218.050 128.115 218.065 ;
        RECT 129.110 218.050 129.410 224.760 ;
        RECT 127.785 217.750 129.410 218.050 ;
        RECT 127.785 217.735 128.115 217.750 ;
        RECT 125.415 211.185 125.745 211.515 ;
        RECT 132.790 210.115 133.090 224.760 ;
        RECT 132.775 209.785 133.105 210.115 ;
        RECT 136.470 209.215 136.770 224.760 ;
        RECT 136.455 208.885 136.785 209.215 ;
        RECT 140.150 208.315 140.450 224.760 ;
        RECT 140.135 207.985 140.465 208.315 ;
        RECT 143.830 207.515 144.130 224.760 ;
        RECT 143.815 207.185 144.145 207.515 ;
        RECT 147.510 206.865 147.810 224.760 ;
        RECT 147.495 206.535 147.825 206.865 ;
        RECT 105.745 160.250 107.255 160.255 ;
        RECT 105.745 158.750 134.750 160.250 ;
        RECT 105.745 158.745 107.255 158.750 ;
        RECT 133.250 152.500 134.750 158.750 ;
        RECT 133.000 150.000 135.000 152.500 ;
        RECT 155.250 44.695 157.150 44.850 ;
        RECT 155.245 44.500 157.150 44.695 ;
        RECT 155.245 44.095 157.160 44.500 ;
        RECT 102.170 37.970 103.230 39.030 ;
        RECT 100.620 36.470 101.680 37.530 ;
        RECT 89.900 1.000 90.920 3.500 ;
        RECT 112.400 1.000 113.000 4.050 ;
        RECT 134.480 1.000 135.080 7.000 ;
        RECT 155.250 6.450 157.160 44.095 ;
        RECT 156.500 1.400 157.160 6.450 ;
        RECT 156.560 1.000 157.160 1.400 ;
        RECT 89.900 0.800 90.320 1.000 ;
  END
END tt_um_emilian_rf_playground
END LIBRARY

