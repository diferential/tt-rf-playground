magic
tech sky130A
magscale 1 2
timestamp 1717256045
<< locali >>
rect -1420 1180 2440 1240
rect -260 940 -200 1180
rect 1200 940 1280 1180
rect -260 660 -200 820
rect 1200 660 1280 820
rect -1420 600 2440 660
rect -150 -310 -60 120
rect 2100 -310 2190 110
<< viali >>
rect 750 1000 800 1050
rect -575 863 -541 897
rect -380 860 -320 920
rect -50 850 0 900
rect 340 850 390 900
rect 560 860 610 910
rect 870 860 920 910
rect 1060 860 1140 900
rect -140 300 -60 380
rect 2120 320 2200 400
rect 18 163 52 197
rect 102 113 148 263
rect 288 163 322 197
rect 372 113 418 263
rect 558 163 592 197
rect 642 113 688 263
rect 828 163 862 197
rect 912 113 958 263
rect 1098 163 1132 197
rect 1182 113 1228 263
rect 1368 163 1402 197
rect 1452 113 1498 263
rect 1638 163 1672 197
rect 1722 113 1768 263
rect 1908 163 1942 197
rect 1992 113 2038 263
rect -140 -540 -60 -460
rect 0 -463 46 -313
rect 96 -397 130 -363
rect 270 -463 316 -313
rect 366 -397 400 -363
rect 540 -463 586 -313
rect 636 -397 670 -363
rect 810 -463 856 -313
rect 906 -397 940 -363
rect 1080 -463 1126 -313
rect 1176 -397 1210 -363
rect 1350 -463 1396 -313
rect 1446 -397 1480 -363
rect 1620 -463 1666 -313
rect 1716 -397 1750 -363
rect 1890 -463 1936 -313
rect 1986 -397 2020 -363
rect 2120 -540 2200 -460
<< metal1 >>
rect -2100 1220 2250 1240
rect -2100 1160 -1300 1220
rect -1210 1160 2250 1220
rect -2100 1150 2250 1160
rect 2380 1150 2440 1240
rect -2100 1140 2440 1150
rect -2100 1000 -320 1080
rect -400 926 -320 1000
rect -50 1056 810 1060
rect -50 1050 812 1056
rect -50 1010 750 1050
rect -400 920 -308 926
rect -2100 910 -480 920
rect -2100 897 -470 910
rect -2100 863 -575 897
rect -541 863 -470 897
rect -2100 840 -470 863
rect -400 860 -380 920
rect -320 860 -308 920
rect -50 906 0 1010
rect 738 1000 750 1010
rect 800 1000 812 1050
rect 738 994 812 1000
rect 1060 920 1160 940
rect 548 910 622 916
rect 858 910 932 916
rect 340 906 390 910
rect -392 854 -308 860
rect -62 900 12 906
rect -62 850 -50 900
rect 0 850 12 900
rect -62 844 12 850
rect 328 900 402 906
rect 328 850 340 900
rect 390 850 402 900
rect 548 860 560 910
rect 610 860 870 910
rect 920 860 932 910
rect 1060 906 1080 920
rect 548 854 622 860
rect 858 854 932 860
rect 1048 900 1080 906
rect 1048 860 1060 900
rect 1140 860 1160 920
rect 1048 854 1160 860
rect 328 844 402 850
rect -520 810 -470 840
rect 340 810 390 844
rect 1060 840 1160 854
rect -520 760 390 810
rect -2100 680 2440 700
rect -2100 620 -1130 680
rect -1030 620 -940 680
rect -840 620 2440 680
rect -2100 600 2440 620
rect -2100 440 -1900 600
rect -1300 520 2220 540
rect -1300 440 -500 520
rect -510 420 -500 440
rect -220 440 2220 520
rect -220 420 -210 440
rect 2108 400 2212 406
rect -1296 330 -1290 390
rect -1230 380 -1224 390
rect -140 386 -60 400
rect -152 380 -48 386
rect 2108 380 2120 400
rect -1230 330 -140 380
rect -1290 320 -140 330
rect -152 300 -140 320
rect -60 320 2120 380
rect 2200 320 2212 400
rect -60 300 -48 320
rect 2108 314 2212 320
rect -152 294 -48 300
rect -140 260 -60 294
rect 96 263 154 275
rect -2100 120 -1340 260
rect -1260 120 -1240 260
rect -60 203 60 220
rect -60 200 64 203
rect -60 140 -40 200
rect 20 197 64 200
rect 52 163 64 197
rect 20 157 64 163
rect 20 140 60 157
rect 96 113 102 263
rect 148 210 154 263
rect 366 263 424 275
rect 148 203 330 210
rect 148 197 334 203
rect 148 163 288 197
rect 322 163 334 197
rect 148 157 334 163
rect 148 150 330 157
rect 148 113 154 150
rect 96 101 154 113
rect 366 113 372 263
rect 418 210 424 263
rect 636 263 694 275
rect 418 203 600 210
rect 418 197 604 203
rect 418 163 558 197
rect 592 163 604 197
rect 418 157 604 163
rect 418 150 600 157
rect 418 113 424 150
rect 366 101 424 113
rect 636 113 642 263
rect 688 210 694 263
rect 906 263 964 275
rect 688 203 870 210
rect 688 197 874 203
rect 688 163 828 197
rect 862 163 874 197
rect 688 157 874 163
rect 688 150 870 157
rect 688 113 694 150
rect 636 101 694 113
rect 906 113 912 263
rect 958 210 964 263
rect 1176 263 1234 275
rect 958 203 1140 210
rect 958 200 1144 203
rect 1060 197 1144 200
rect 1060 163 1098 197
rect 1132 163 1144 197
rect 1060 157 1144 163
rect 1060 150 1140 157
rect 1060 140 1070 150
rect 958 113 964 140
rect 906 101 964 113
rect 1176 113 1182 263
rect 1228 210 1234 263
rect 1446 263 1504 275
rect 1228 203 1410 210
rect 1228 197 1414 203
rect 1228 163 1368 197
rect 1402 163 1414 197
rect 1228 157 1414 163
rect 1228 150 1410 157
rect 1228 113 1234 150
rect 1176 101 1234 113
rect 1446 113 1452 263
rect 1498 210 1504 263
rect 1716 263 1774 275
rect 1498 203 1680 210
rect 1498 197 1684 203
rect 1498 163 1638 197
rect 1672 163 1684 197
rect 1498 157 1684 163
rect 1498 150 1680 157
rect 1498 113 1504 150
rect 1446 101 1504 113
rect 1716 113 1722 263
rect 1768 210 1774 263
rect 1986 263 2044 275
rect 1768 203 1950 210
rect 1768 197 1954 203
rect 1768 163 1908 197
rect 1942 163 1954 197
rect 1768 157 1954 163
rect 1768 150 1950 157
rect 1768 113 1774 150
rect 1716 101 1774 113
rect 1986 113 1992 263
rect 2038 230 2044 263
rect 2120 260 2200 314
rect 2038 220 2090 230
rect 2070 160 2090 220
rect 2038 150 2090 160
rect 2038 113 2044 150
rect 1986 101 2044 113
rect -1300 -140 -1140 0
rect -1000 -40 2220 0
rect -1000 -140 -940 -40
rect -840 -140 2220 -40
rect -1300 -200 2220 -140
rect -6 -313 52 -301
rect -6 -340 0 -313
rect -50 -400 -40 -340
rect -50 -420 0 -400
rect -152 -460 -48 -454
rect -1290 -470 -1230 -464
rect -152 -470 -140 -460
rect -1230 -530 -140 -470
rect -1290 -536 -1230 -530
rect -152 -540 -140 -530
rect -60 -520 -48 -460
rect -6 -463 0 -420
rect 46 -463 52 -313
rect 264 -313 322 -301
rect 264 -350 270 -313
rect 90 -357 270 -350
rect 84 -363 270 -357
rect 84 -397 96 -363
rect 130 -397 270 -363
rect 84 -403 270 -397
rect 90 -410 270 -403
rect -6 -475 52 -463
rect 264 -463 270 -410
rect 316 -463 322 -313
rect 534 -313 592 -301
rect 534 -350 540 -313
rect 360 -357 540 -350
rect 354 -363 540 -357
rect 354 -397 366 -363
rect 400 -397 540 -363
rect 354 -403 540 -397
rect 360 -410 540 -403
rect 264 -475 322 -463
rect 534 -463 540 -410
rect 586 -463 592 -313
rect 804 -313 862 -301
rect 804 -350 810 -313
rect 640 -357 810 -350
rect 624 -363 810 -357
rect 624 -397 636 -363
rect 670 -397 810 -363
rect 624 -403 810 -397
rect 640 -410 810 -403
rect 534 -475 592 -463
rect 804 -463 810 -410
rect 856 -463 862 -313
rect 1074 -313 1132 -301
rect 1074 -350 1080 -313
rect 900 -357 1080 -350
rect 894 -363 1080 -357
rect 894 -397 906 -363
rect 940 -397 1080 -363
rect 894 -403 1080 -397
rect 900 -410 1080 -403
rect 804 -475 862 -463
rect 1074 -463 1080 -410
rect 1126 -463 1132 -313
rect 1344 -313 1402 -301
rect 1344 -350 1350 -313
rect 1170 -357 1350 -350
rect 1164 -363 1350 -357
rect 1164 -397 1176 -363
rect 1210 -397 1350 -363
rect 1164 -403 1350 -397
rect 1170 -410 1350 -403
rect 1074 -475 1132 -463
rect 1344 -463 1350 -410
rect 1396 -463 1402 -313
rect 1614 -313 1672 -301
rect 1614 -350 1620 -313
rect 1440 -357 1620 -350
rect 1434 -363 1620 -357
rect 1434 -397 1446 -363
rect 1480 -397 1620 -363
rect 1434 -403 1620 -397
rect 1440 -410 1620 -403
rect 1344 -475 1402 -463
rect 1614 -463 1620 -410
rect 1666 -463 1672 -313
rect 1884 -313 1942 -301
rect 1884 -350 1890 -313
rect 1710 -357 1890 -350
rect 1704 -363 1890 -357
rect 1704 -397 1716 -363
rect 1750 -397 1890 -363
rect 1704 -403 1890 -397
rect 1710 -410 1890 -403
rect 1614 -475 1672 -463
rect 1884 -463 1890 -410
rect 1936 -463 1942 -313
rect 1970 -350 2080 -340
rect 1970 -363 2010 -350
rect 1970 -397 1986 -363
rect 1970 -410 2010 -397
rect 2070 -410 2080 -350
rect 1970 -420 2080 -410
rect 1884 -475 1942 -463
rect 2108 -460 2212 -454
rect 2108 -520 2120 -460
rect -60 -540 2120 -520
rect 2200 -540 2212 -460
rect -152 -546 2120 -540
rect -140 -580 2120 -546
rect 2180 -546 2212 -540
rect 2180 -580 2200 -546
rect -510 -600 -500 -580
rect -2120 -680 -500 -600
rect -220 -640 -210 -580
rect -140 -600 -60 -580
rect 2120 -600 2200 -580
rect -220 -680 2220 -640
rect -2120 -740 2220 -680
<< via1 >>
rect -1300 1160 -1210 1220
rect 2250 1150 2380 1240
rect 1080 900 1140 920
rect 1080 860 1140 900
rect -1130 620 -1030 680
rect -940 620 -840 680
rect -500 420 -220 520
rect -1290 330 -1230 390
rect 2120 330 2180 390
rect -1340 120 -1260 260
rect -40 197 20 200
rect -40 163 18 197
rect 18 163 20 197
rect -40 140 20 163
rect 940 140 958 200
rect 958 140 1060 200
rect 2010 160 2038 220
rect 2038 160 2070 220
rect -1140 -140 -1000 0
rect -940 -140 -840 -40
rect -40 -400 0 -340
rect 0 -400 20 -340
rect -1290 -530 -1230 -470
rect 2010 -363 2070 -350
rect 2010 -397 2020 -363
rect 2020 -397 2070 -363
rect 2010 -410 2070 -397
rect 2120 -540 2180 -520
rect 2120 -580 2180 -540
rect -500 -680 -220 -580
<< metal2 >>
rect 2250 1240 2380 1250
rect -1340 1230 -1230 1240
rect -1340 1220 -1210 1230
rect -1340 1160 -1300 1220
rect -1340 1150 -1210 1160
rect -1340 390 -1230 1150
rect 2250 1140 2380 1150
rect 1060 920 1140 940
rect 1060 860 1080 920
rect 1060 840 1140 860
rect -1340 330 -1290 390
rect -1340 260 -1230 330
rect -1260 120 -1230 260
rect -1340 110 -1230 120
rect -1290 -470 -1230 110
rect -1170 680 -800 700
rect -1170 620 -1130 680
rect -1030 620 -940 680
rect -840 620 -800 680
rect -1170 0 -800 620
rect -1170 -140 -1140 0
rect -1000 -40 -800 0
rect -1000 -140 -940 -40
rect -840 -140 -800 -40
rect -1170 -190 -800 -140
rect -500 520 -220 540
rect -1296 -530 -1290 -470
rect -1230 -530 -1224 -470
rect -500 -580 -220 420
rect 1080 220 1140 840
rect 2280 400 2350 1140
rect 2120 390 2350 400
rect 2180 330 2350 390
rect 2120 320 2350 330
rect 2120 310 2180 320
rect 2010 220 2070 230
rect -50 200 30 220
rect -50 140 -40 200
rect 20 140 30 200
rect 900 200 1140 220
rect 900 140 940 200
rect 1060 140 1140 200
rect 2000 160 2010 220
rect 2070 160 2080 220
rect 2000 150 2080 160
rect -40 -340 20 140
rect 940 130 1060 140
rect 2000 110 2070 150
rect 2010 -340 2070 110
rect -50 -400 -40 -340
rect 20 -400 30 -340
rect -50 -420 30 -400
rect 2000 -350 2080 -340
rect 2000 -410 2010 -350
rect 2070 -410 2080 -350
rect 2000 -420 2080 -410
rect 2120 -500 2180 -490
rect 2280 -500 2350 320
rect 2120 -520 2350 -500
rect 2114 -580 2120 -520
rect 2180 -580 2350 -520
rect -500 -720 -220 -680
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 -198 0 -1 -148
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_1
timestamp 1707688321
transform 1 0 -1302 0 1 -52
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 878 0 1 648
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 458 0 1 648
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 -142 0 1 648
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 -962 0 1 648
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1338 0 1 648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1707688321
transform 1 0 -2102 0 1 648
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1828 0 1 -52
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1707688321
transform 1 0 -62 0 1 -52
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1707688321
transform 1 0 208 0 1 -52
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1707688321
transform 1 0 478 0 1 -52
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1707688321
transform 1 0 748 0 1 -52
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1707688321
transform 1 0 1018 0 1 -52
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1707688321
transform 1 0 1288 0 1 -52
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1707688321
transform 1 0 1558 0 1 -52
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1707688321
transform -1 0 1560 0 -1 -148
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1707688321
transform -1 0 2100 0 -1 -148
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1707688321
transform -1 0 1830 0 -1 -148
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_11
timestamp 1707688321
transform -1 0 750 0 -1 -148
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_12
timestamp 1707688321
transform -1 0 1290 0 -1 -148
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_13
timestamp 1707688321
transform -1 0 1020 0 -1 -148
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_14
timestamp 1707688321
transform -1 0 210 0 -1 -148
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_15
timestamp 1707688321
transform -1 0 480 0 -1 -148
box -38 -48 314 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 -60 0 -1 -148
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_1
timestamp 1707688321
transform 1 0 2098 0 1 -52
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_2
timestamp 1707688321
transform 1 0 -142 0 1 -52
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_3
timestamp 1707688321
transform -1 0 2190 0 -1 -148
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_4
timestamp 1707688321
transform 1 0 -272 0 1 648
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_5
timestamp 1707688321
transform 1 0 1198 0 1 648
box -38 -48 130 592
<< labels >>
flabel metal1 -2120 -740 -1980 -600 0 FreeSans 1600 0 0 0 VIN
port 0 nsew
flabel metal1 -2100 1000 -2000 1080 0 FreeSans 1600 0 0 0 VOUT
port 1 nsew
flabel metal1 -2100 840 -2000 920 0 FreeSans 1600 0 0 0 VOUT_N
port 2 nsew
flabel metal1 -2100 120 -1960 260 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal1 -2100 440 -1960 580 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
<< end >>
