magic
tech sky130A
magscale 1 2
timestamp 1717254928
<< nwell >>
rect -480 -1060 -380 500
rect -980 -1140 -380 -1060
rect -980 -1160 -420 -1140
<< locali >>
rect -1400 3180 -700 3200
rect -1400 2760 10520 3180
rect -1400 2620 -280 2760
rect -1400 2600 -220 2620
rect -1400 2460 100 2600
rect -1400 1920 -760 2460
rect -380 1920 100 2460
rect 9600 2500 10200 2600
rect 9600 2300 9900 2400
rect -1400 1220 100 1920
rect -1400 1120 -380 1220
rect -200 1200 100 1220
rect -1400 880 -900 1120
rect -1400 260 -800 880
rect -1400 -80 -900 260
rect -680 200 -540 980
rect -460 500 -380 1120
rect -1260 -160 -900 -80
rect -1260 -860 -800 -160
rect -1400 -900 -800 -860
rect -1400 -1060 -900 -900
rect -480 -1060 -380 500
rect -1400 -1080 -380 -1060
rect -1400 -1120 -900 -1080
rect -520 -1120 -380 -1080
rect -1400 -1140 -380 -1120
rect -300 1000 0 1100
rect -300 200 -200 1000
rect -100 200 0 1000
rect -300 -300 0 200
rect -300 -1000 -200 -300
rect -100 -1000 0 -300
rect -300 -1100 0 -1000
rect -1400 -1160 -420 -1140
rect -1400 -2300 -900 -1160
rect -300 -1280 -100 -1100
rect -740 -1860 -100 -1280
rect -400 -2300 400 -2251
rect 9800 -2300 9900 2300
rect -1400 -2600 400 -2300
rect 9600 -2400 9900 -2300
rect 10100 -2500 10200 2500
rect 9600 -2600 10200 -2500
rect -1400 -2700 -100 -2600
rect -1400 -3300 10140 -2700
<< viali >>
rect -760 1920 -380 2460
rect 9600 2400 10100 2500
rect -900 -1120 -520 -1080
rect -200 200 -100 1000
rect -200 -1000 -100 -300
rect 9900 -2400 10100 2400
rect 9600 -2500 10100 -2400
<< metal1 >>
rect -1400 3180 -700 3200
rect -1400 2760 10520 3180
rect -1400 2600 -280 2760
rect -1400 2460 0 2600
rect -1400 1920 -760 2460
rect -380 2300 0 2460
rect 9600 2500 10200 2600
rect 9600 2300 9900 2400
rect -380 1920 -200 2300
rect -1400 1300 -200 1920
rect -1400 1220 -300 1300
rect -1400 1140 -380 1220
rect -1400 1120 -820 1140
rect -540 1120 -380 1140
rect -1400 880 -900 1120
rect -740 980 -660 1060
rect -1400 260 -800 880
rect -1400 -80 -900 260
rect -740 200 -540 980
rect -460 500 -380 1120
rect -740 120 -660 200
rect -780 60 -620 120
rect -780 -40 -760 60
rect -660 -40 -620 60
rect -780 -60 -620 -40
rect -740 -80 -660 -60
rect -1260 -160 -900 -80
rect -1260 -860 -800 -160
rect -1400 -900 -800 -860
rect -1400 -1060 -900 -900
rect -760 -980 -660 -80
rect -630 -160 -520 -120
rect -630 -900 -620 -160
rect -540 -900 -520 -160
rect -630 -940 -520 -900
rect -740 -1000 -660 -980
rect -480 -1060 -380 500
rect -1400 -1080 -380 -1060
rect -1400 -1120 -900 -1080
rect -520 -1120 -380 -1080
rect -1400 -1140 -380 -1120
rect -300 1000 0 1100
rect -300 200 -200 1000
rect -100 200 0 1000
rect -300 -300 0 200
rect -300 -1000 -200 -300
rect -100 -1000 0 -300
rect -300 -1100 0 -1000
rect -1400 -1160 -420 -1140
rect -1400 -2300 -900 -1160
rect -300 -1280 -100 -1100
rect -740 -1860 -100 -1280
rect -400 -2300 349 -2251
rect 9800 -2300 9900 2300
rect -1400 -2500 400 -2300
rect 9600 -2400 9900 -2300
rect 10100 -2500 10200 2500
rect -1400 -2549 349 -2500
rect -1400 -2600 200 -2549
rect 9600 -2600 10200 -2500
rect -1400 -2700 -100 -2600
rect -1400 -3300 10140 -2700
<< via1 >>
rect -760 -40 -660 60
rect -620 -900 -540 -160
<< metal2 >>
rect 1800 3090 10530 3190
rect 1800 2565 1900 3090
rect 4200 2890 10330 2990
rect 4200 2585 4300 2890
rect 6600 2690 10090 2790
rect 6600 2600 6700 2690
rect 6580 2585 6720 2600
rect 1796 2475 1805 2565
rect 1895 2475 1904 2565
rect 4196 2495 4205 2585
rect 4295 2495 4304 2585
rect 6580 2495 6605 2585
rect 6695 2495 6720 2585
rect 4200 2490 4300 2495
rect 6580 2480 6720 2495
rect 8980 2570 9120 2600
rect 8980 2565 9930 2570
rect 8980 2475 9005 2565
rect 9095 2475 9930 2565
rect 1800 2470 1900 2475
rect 8980 2470 9930 2475
rect 8980 2460 9120 2470
rect -100 2152 200 2200
rect -1638 1918 200 2152
rect 9679 2140 9761 2161
rect 9400 1980 9761 2140
rect -100 1900 200 1918
rect 2160 1520 2340 1530
rect 2160 1350 2340 1360
rect 4580 1520 4760 1530
rect 4580 1350 4760 1360
rect 6960 1520 7140 1530
rect 6960 1350 7140 1360
rect 9380 1520 9560 1530
rect 9380 1350 9560 1360
rect -820 120 -560 140
rect -300 120 9600 200
rect -820 100 9600 120
rect -820 60 100 100
rect -820 -40 -760 60
rect -660 -40 100 60
rect -820 -80 -560 -40
rect -300 -100 100 -40
rect 300 -100 2200 100
rect 2600 -100 4600 100
rect 5000 -100 7000 100
rect 7400 -100 9300 100
rect 9500 -100 9600 100
rect -620 -160 -540 -150
rect -1400 -780 -620 -180
rect -540 -780 -520 -180
rect -300 -200 9600 -100
rect -620 -910 -540 -900
rect 40 -1340 220 -1330
rect 40 -1510 220 -1500
rect 2460 -1340 2640 -1330
rect 7240 -1340 7420 -1330
rect 2460 -1510 2640 -1500
rect 4840 -1360 5020 -1350
rect 7240 -1510 7420 -1500
rect 4840 -1530 5020 -1520
rect -1400 -1940 -940 -1920
rect -100 -1940 200 -1900
rect -1400 -2014 200 -1940
rect -1638 -2134 200 -2014
rect -1400 -2180 200 -2134
rect 9400 -2034 9576 -1960
rect 9679 -1981 9761 1980
rect 9830 110 9930 2470
rect 9990 310 10090 2690
rect 10230 490 10330 2890
rect 10430 810 10530 3090
rect 10430 710 11376 810
rect 10230 390 11376 490
rect 9990 210 11376 310
rect 9830 10 11376 110
rect 9850 -230 11376 -130
rect 9680 -2034 9760 -1981
rect 9400 -2160 9760 -2034
rect -100 -2200 200 -2180
rect 490 -2510 590 -2501
rect 475 -2610 490 -2515
rect 475 -2920 590 -2610
rect 2890 -2510 2990 -2501
rect 475 -3000 560 -2920
rect 480 -3160 560 -3000
rect 2890 -3010 2990 -2610
rect 5290 -2520 5390 -2510
rect 5290 -2600 5300 -2520
rect 5380 -2600 5390 -2520
rect 5290 -2830 5390 -2600
rect 7660 -2520 7820 -2500
rect 9850 -2510 9950 -230
rect 7660 -2600 7700 -2520
rect 7780 -2600 7820 -2520
rect 7660 -2610 7820 -2600
rect 9690 -2610 9950 -2510
rect 7660 -2710 9950 -2610
rect 10050 -430 11376 -330
rect 7660 -2720 7820 -2710
rect 10050 -2830 10150 -430
rect 10290 -630 11376 -530
rect 10290 -1160 10390 -630
rect 10450 -850 11376 -750
rect 10450 -1160 10550 -850
rect 10288 -1840 10392 -1160
rect 10450 -1840 10552 -1160
rect 5290 -2930 10150 -2830
rect 10290 -3010 10390 -1840
rect 2880 -3110 10390 -3010
rect 480 -3210 565 -3160
rect 10450 -3210 10550 -1840
rect 480 -3300 10550 -3210
<< via2 >>
rect 1805 2475 1895 2565
rect 4205 2495 4295 2585
rect 6605 2495 6695 2585
rect 9005 2475 9095 2565
rect 2160 1360 2340 1520
rect 4580 1360 4760 1520
rect 6960 1360 7140 1520
rect 9380 1360 9560 1520
rect 100 -100 300 100
rect 2200 -100 2600 100
rect 4600 -100 5000 100
rect 7000 -100 7400 100
rect 9300 -100 9500 100
rect 40 -1500 220 -1340
rect 2460 -1500 2640 -1340
rect 4840 -1520 5020 -1360
rect 7240 -1500 7420 -1340
rect 490 -2610 590 -2510
rect 2890 -2610 2990 -2510
rect 5300 -2600 5380 -2520
rect 7700 -2600 7780 -2520
<< metal3 >>
rect 4200 2585 4300 2590
rect 1800 2565 1900 2570
rect 1800 2475 1805 2565
rect 1895 2475 1900 2565
rect 4200 2495 4205 2585
rect 4295 2495 4300 2585
rect 4200 2490 4300 2495
rect 6600 2585 6700 2590
rect 6600 2495 6605 2585
rect 6695 2495 6700 2585
rect 6600 2490 6700 2495
rect 9000 2565 9100 2570
rect 1800 2470 1900 2475
rect 9000 2475 9005 2565
rect 9095 2475 9100 2565
rect 9000 2470 9100 2475
rect 2100 1520 2400 1600
rect 2100 1360 2160 1520
rect 2340 1360 2400 1520
rect 2100 200 2400 1360
rect 4500 1520 4800 1600
rect 4500 1360 4580 1520
rect 4760 1360 4800 1520
rect 4500 200 4800 1360
rect 6900 1520 7200 1600
rect 6900 1360 6960 1520
rect 7140 1360 7200 1520
rect 6900 200 7200 1360
rect 9300 1520 9600 1600
rect 9300 1360 9380 1520
rect 9560 1360 9600 1520
rect 9300 200 9600 1360
rect 0 100 400 200
rect 0 -100 100 100
rect 300 -100 400 100
rect 0 -200 400 -100
rect 2100 100 2700 200
rect 2100 -100 2200 100
rect 2600 -100 2700 100
rect 2100 -200 2700 -100
rect 4500 100 5100 200
rect 4500 -100 4600 100
rect 5000 -100 5100 100
rect 4500 -200 5100 -100
rect 6900 100 7500 200
rect 6900 -100 7000 100
rect 7400 -100 7500 100
rect 6900 -200 7500 -100
rect 9200 100 9600 200
rect 9200 -100 9300 100
rect 9500 -100 9600 100
rect 9200 -200 9600 -100
rect 0 -1340 300 -200
rect 0 -1500 40 -1340
rect 220 -1500 300 -1340
rect 0 -1600 300 -1500
rect 2400 -1340 2700 -200
rect 2400 -1500 2460 -1340
rect 2640 -1500 2700 -1340
rect 2400 -1600 2700 -1500
rect 4800 -1360 5100 -200
rect 4800 -1520 4840 -1360
rect 5020 -1520 5100 -1360
rect 4800 -1600 5100 -1520
rect 7200 -1340 7500 -200
rect 7200 -1500 7240 -1340
rect 7420 -1500 7500 -1340
rect 7200 -1600 7500 -1500
rect 485 -2510 595 -2505
rect 485 -2610 490 -2510
rect 590 -2610 595 -2510
rect 485 -2615 595 -2610
rect 2885 -2510 2995 -2505
rect 2885 -2610 2890 -2510
rect 2990 -2610 2995 -2510
rect 5290 -2520 5390 -2515
rect 5290 -2600 5300 -2520
rect 5380 -2600 5390 -2520
rect 5290 -2605 5390 -2600
rect 7690 -2520 7790 -2515
rect 7690 -2600 7700 -2520
rect 7780 -2600 7790 -2520
rect 7690 -2605 7790 -2600
rect 2885 -2615 2995 -2610
use idac1cell  idac1cell_0
timestamp 1713553032
transform -1 0 2000 0 -1 200
box -400 200 2000 2800
use idac1cell  idac1cell_1
timestamp 1713553032
transform 1 0 400 0 1 -200
box -400 200 2000 2800
use idac1cell  idac1cell_2
timestamp 1713553032
transform 1 0 2800 0 1 -200
box -400 200 2000 2800
use idac1cell  idac1cell_3
timestamp 1713553032
transform 1 0 5200 0 1 -200
box -400 200 2000 2800
use idac1cell  idac1cell_4
timestamp 1713553032
transform 1 0 7600 0 1 -200
box -400 200 2000 2800
use idac1cell  idac1cell_5
timestamp 1713553032
transform -1 0 9200 0 -1 200
box -400 200 2000 2800
use idac1cell  idac1cell_6
timestamp 1713553032
transform -1 0 6800 0 -1 200
box -400 200 2000 2800
use idac1cell  idac1cell_7
timestamp 1713553032
transform -1 0 4400 0 -1 200
box -400 200 2000 2800
use sky130_fd_pr__pfet_01v8_lvt_ZJ8M88  sky130_fd_pr__pfet_01v8_lvt_ZJ8M88_0
timestamp 1713499374
transform 1 0 -694 0 1 -531
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_lvt_ZJ82X3  sky130_fd_pr__pfet_01v8_lvt_ZJ82X3_0
timestamp 1713499374
transform 1 0 -694 0 1 579
box -296 -619 296 619
<< labels >>
flabel metal2 -100 1900 200 2200 0 FreeSans 1600 0 0 0 VREF_IN
port 8 nsew
flabel metal2 10520 720 10600 800 0 FreeSans 1600 0 0 0 VCMD0
port 0 nsew
flabel metal2 10520 400 10600 480 0 FreeSans 1600 0 0 0 VCMD1
port 1 nsew
flabel metal2 10520 220 10600 300 0 FreeSans 1600 0 0 0 VCMD2
port 2 nsew
flabel metal2 10520 20 10600 100 0 FreeSans 1600 0 0 0 VCMD3
port 3 nsew
flabel metal2 10520 -220 10600 -140 0 FreeSans 1600 0 0 0 VCMD4
port 4 nsew
flabel metal2 10520 -420 10600 -340 0 FreeSans 1600 0 0 0 VCMD5
port 5 nsew
flabel metal2 10520 -620 10600 -540 0 FreeSans 1600 0 0 0 VCMD6
port 6 nsew
flabel metal2 10540 -840 10620 -760 0 FreeSans 1600 0 0 0 VCMD7
port 7 nsew
flabel metal2 -1400 -780 -1280 -180 0 FreeSans 1600 0 0 0 IOUT_P
port 10 nsew
flabel metal2 -1340 -2120 -1020 -1960 0 FreeSans 1600 0 0 0 VREF_OUT
port 9 nsew
flabel metal1 -1314 2702 -664 3086 0 FreeSans 1600 0 0 0 VDD
port 11 nsew
<< end >>
