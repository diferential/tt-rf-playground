magic
tech sky130A
timestamp 1719784978
<< pwell >>
rect 0 0 360 170
<< nmos >>
rect 40 50 55 95
rect 95 50 110 95
rect 135 50 150 95
rect 190 50 205 95
rect 230 50 245 95
rect 285 50 300 95
<< ndiff >>
rect 5 85 40 95
rect 5 65 10 85
rect 30 65 40 85
rect 5 50 40 65
rect 55 85 95 95
rect 55 65 65 85
rect 85 65 95 85
rect 55 50 95 65
rect 110 50 135 95
rect 150 85 190 95
rect 150 65 160 85
rect 180 65 190 85
rect 150 50 190 65
rect 205 50 230 95
rect 245 80 285 95
rect 245 60 255 80
rect 275 60 285 80
rect 245 50 285 60
rect 300 80 335 95
rect 300 60 310 80
rect 330 60 335 80
rect 300 50 335 60
<< ndiffc >>
rect 10 65 30 85
rect 65 65 85 85
rect 160 65 180 85
rect 255 60 275 80
rect 310 60 330 80
<< poly >>
rect 40 95 55 170
rect 95 95 110 170
rect 175 140 205 150
rect 175 120 180 140
rect 200 120 205 140
rect 175 110 205 120
rect 135 95 150 110
rect 190 95 205 110
rect 230 95 245 170
rect 285 95 300 170
rect 40 0 55 50
rect 95 0 110 50
rect 135 40 150 50
rect 135 30 165 40
rect 190 35 205 50
rect 135 10 140 30
rect 160 10 165 30
rect 135 0 165 10
rect 230 0 245 50
rect 285 0 300 50
<< polycont >>
rect 180 120 200 140
rect 140 10 160 30
<< locali >>
rect 0 140 210 150
rect 0 120 180 140
rect 200 120 210 140
rect 0 115 210 120
rect 0 85 40 115
rect 0 65 10 85
rect 30 65 40 85
rect 0 0 40 65
rect 60 85 90 95
rect 60 65 65 85
rect 85 65 90 85
rect 60 50 90 65
rect 155 85 185 95
rect 155 65 160 85
rect 180 65 185 85
rect 155 50 185 65
rect 250 80 280 95
rect 250 60 255 80
rect 275 60 280 80
rect 250 50 280 60
rect 300 80 340 150
rect 300 60 310 80
rect 330 60 340 80
rect 300 30 340 60
rect 130 10 140 30
rect 160 10 340 30
rect 130 0 340 10
<< viali >>
rect 10 65 30 85
rect 65 65 85 85
rect 160 65 180 85
rect 255 60 275 80
rect 310 60 330 80
<< metal1 >>
rect 0 105 360 120
rect 0 85 40 90
rect 65 88 85 105
rect 0 65 10 85
rect 30 65 40 85
rect 0 60 40 65
rect 59 85 91 88
rect 59 65 65 85
rect 85 65 91 85
rect 59 62 91 65
rect 150 60 155 90
rect 185 60 190 90
rect 249 80 281 83
rect 249 60 255 80
rect 275 60 281 80
rect 249 57 281 60
rect 300 80 340 85
rect 300 60 310 80
rect 330 60 340 80
rect 255 40 275 57
rect 300 55 340 60
rect 0 25 360 40
<< via1 >>
rect 155 85 185 90
rect 155 65 160 85
rect 160 65 180 85
rect 180 65 185 85
rect 155 60 185 65
<< metal2 >>
rect 155 90 185 170
rect 155 0 185 60
<< labels >>
flabel ndiffc 160 65 180 85 0 FreeSans 80 90 0 0 VS
flabel ndiff 70 65 90 85 0 FreeSans 80 90 0 0 BL
flabel ndiff 255 65 275 85 0 FreeSans 80 90 0 0 BLB
flabel poly 230 145 245 160 0 FreeSans 80 90 0 0 RDB
flabel poly 95 10 110 25 0 FreeSans 80 90 0 0 RD
flabel poly 285 145 300 160 0 FreeSans 80 90 0 0 WR
flabel poly 40 10 55 25 0 FreeSans 80 90 0 0 WRB
flabel locali 0 130 15 145 0 FreeSans 80 90 0 0 VGB
flabel locali 325 10 340 25 0 FreeSans 80 90 0 0 VG
<< properties >>
string FIXED_BBOX 0 0 360 170
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
