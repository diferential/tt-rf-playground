magic
tech sky130A
magscale 1 2
timestamp 1723170491
<< pwell >>
rect -140 -400 2710 400
<< psubdiff >>
rect -120 340 470 380
rect 2140 340 2680 380
rect -120 -340 -80 340
rect 2640 -340 2680 340
rect -120 -380 450 -340
rect 2120 -380 2680 -340
<< psubdiffcont >>
rect 470 340 2140 380
rect 450 -380 2120 -340
<< locali >>
rect -120 340 470 380
rect 2140 340 2680 380
rect -120 -340 -80 340
rect 140 -170 180 120
rect 380 -170 420 120
rect 620 -170 660 120
rect 860 -170 900 120
rect 1100 -170 1140 120
rect 1340 -170 1380 120
rect 1580 -170 1620 120
rect 1820 -170 1860 120
rect 2060 -170 2100 120
rect 2300 -170 2340 120
rect 2540 -170 2580 120
rect 2640 -340 2680 340
rect -120 -370 410 -340
rect -120 -380 450 -370
rect 2120 -380 2680 -340
<< viali >>
rect 410 -340 510 -290
rect 1130 -340 1230 -290
rect 1370 -340 1470 -290
rect 410 -370 450 -340
rect 450 -370 510 -340
rect 1130 -370 1230 -340
rect 1370 -370 1470 -340
<< metal1 >>
rect 670 310 680 320
rect -20 270 680 310
rect -20 30 20 270
rect 50 160 60 220
rect 120 160 130 220
rect 220 30 260 270
rect 290 160 300 220
rect 360 160 370 220
rect 460 30 500 270
rect 670 260 680 270
rect 740 260 750 320
rect 1170 310 1230 490
rect 940 270 1460 310
rect 530 160 540 220
rect 600 160 610 220
rect 700 30 740 260
rect 770 160 780 220
rect 840 160 850 220
rect 940 30 980 270
rect 1170 260 1230 270
rect 1010 160 1020 220
rect 1080 160 1090 220
rect 1180 30 1220 260
rect 1250 160 1260 220
rect 1320 160 1330 220
rect 1420 30 1460 270
rect 1510 220 1570 480
rect 1640 260 1650 320
rect 1710 310 1720 320
rect 1710 270 2420 310
rect 1710 260 1720 270
rect 1490 160 1500 220
rect 1560 160 1570 220
rect 1660 30 1700 260
rect 1730 160 1740 220
rect 1800 160 1810 220
rect 1900 30 1940 270
rect 1970 160 1980 220
rect 2040 160 2050 220
rect 2140 30 2180 270
rect 2210 160 2220 220
rect 2280 160 2290 220
rect 2380 30 2420 270
rect 2450 160 2460 220
rect 2520 160 2530 220
rect -20 -290 20 -80
rect -50 -350 -40 -290
rect 20 -350 30 -290
rect -20 -380 20 -350
rect 70 -910 110 -210
rect 220 -290 260 -80
rect 190 -350 200 -290
rect 260 -350 270 -290
rect 220 -380 260 -350
rect 310 -910 350 -210
rect 460 -284 500 -80
rect 398 -290 522 -284
rect 398 -370 410 -290
rect 510 -370 522 -290
rect 398 -376 522 -370
rect 460 -380 500 -376
rect 550 -790 590 -210
rect 700 -290 740 -80
rect 670 -350 680 -290
rect 740 -350 750 -290
rect 700 -380 740 -350
rect 790 -670 830 -210
rect 940 -290 980 -80
rect 910 -350 920 -290
rect 980 -350 990 -290
rect 940 -380 980 -350
rect 1030 -430 1070 -210
rect 1180 -284 1220 -80
rect 1118 -290 1242 -284
rect 1118 -370 1130 -290
rect 1230 -370 1242 -290
rect 1118 -376 1242 -370
rect 1180 -380 1220 -376
rect 1010 -490 1020 -430
rect 1080 -490 1090 -430
rect 770 -730 780 -670
rect 840 -730 850 -670
rect 530 -850 540 -790
rect 600 -850 610 -790
rect 50 -970 60 -910
rect 120 -970 130 -910
rect 290 -970 300 -910
rect 360 -970 370 -910
rect 550 -970 590 -850
rect 790 -970 830 -730
rect 1030 -970 1070 -490
rect 1270 -550 1310 -210
rect 1420 -284 1460 -80
rect 1358 -290 1482 -284
rect 1358 -370 1370 -290
rect 1470 -370 1482 -290
rect 1358 -376 1482 -370
rect 1420 -380 1460 -376
rect 1510 -550 1550 -210
rect 1660 -290 1700 -80
rect 1630 -350 1640 -290
rect 1700 -350 1710 -290
rect 1660 -380 1700 -350
rect 1750 -430 1790 -210
rect 1900 -290 1940 -80
rect 1870 -350 1880 -290
rect 1940 -350 1950 -290
rect 1900 -380 1940 -350
rect 1730 -490 1740 -430
rect 1800 -490 1810 -430
rect 1250 -610 1260 -550
rect 1320 -610 1330 -550
rect 1490 -610 1500 -550
rect 1560 -610 1570 -550
rect 1270 -970 1310 -610
rect 1510 -970 1550 -610
rect 1750 -970 1790 -490
rect 1990 -790 2030 -210
rect 2140 -290 2180 -80
rect 2110 -350 2120 -290
rect 2180 -350 2190 -290
rect 2140 -380 2180 -350
rect 1970 -850 1980 -790
rect 2040 -850 2050 -790
rect 1990 -970 2030 -850
rect 2230 -910 2270 -210
rect 2380 -290 2420 -80
rect 2350 -350 2360 -290
rect 2420 -350 2430 -290
rect 2380 -380 2420 -350
rect 2470 -910 2510 -210
rect 2210 -970 2220 -910
rect 2280 -970 2290 -910
rect 2450 -970 2460 -910
rect 2520 -970 2530 -910
<< via1 >>
rect 60 160 120 220
rect 300 160 360 220
rect 680 260 740 320
rect 540 160 600 220
rect 780 160 840 220
rect 1020 160 1080 220
rect 1260 160 1320 220
rect 1650 260 1710 320
rect 1500 160 1560 220
rect 1740 160 1800 220
rect 1980 160 2040 220
rect 2220 160 2280 220
rect 2460 160 2520 220
rect -40 -350 20 -290
rect 200 -350 260 -290
rect 440 -350 500 -290
rect 680 -350 740 -290
rect 920 -350 980 -290
rect 1160 -350 1220 -290
rect 1020 -490 1080 -430
rect 780 -730 840 -670
rect 540 -850 600 -790
rect 60 -970 120 -910
rect 300 -970 360 -910
rect 1400 -350 1460 -290
rect 1640 -350 1700 -290
rect 1880 -350 1940 -290
rect 1740 -490 1800 -430
rect 1260 -610 1320 -550
rect 1500 -610 1560 -550
rect 2120 -350 2180 -290
rect 1980 -850 2040 -790
rect 2360 -350 2420 -290
rect 2220 -970 2280 -910
rect 2460 -970 2520 -910
<< metal2 >>
rect 680 320 740 330
rect 940 320 1000 490
rect 1650 320 1710 330
rect 740 260 1650 320
rect 680 250 740 260
rect 1650 250 1710 260
rect 60 220 120 230
rect -20 160 60 200
rect 300 220 360 230
rect 120 160 300 200
rect 540 220 600 230
rect 360 160 540 200
rect 780 220 840 230
rect 600 160 780 200
rect 1020 220 1080 230
rect 840 160 1020 200
rect 1260 220 1320 230
rect 1080 160 1260 200
rect 1500 220 1560 230
rect 1320 160 1500 200
rect 1740 220 1800 230
rect 1560 160 1740 200
rect 1980 220 2040 230
rect 1800 160 1980 200
rect 2220 220 2280 230
rect 2040 160 2220 200
rect 2460 220 2520 230
rect 2280 160 2460 200
rect 2520 160 2580 200
rect -20 150 2580 160
rect -40 -290 20 -280
rect 200 -290 260 -280
rect 440 -290 500 -280
rect 680 -290 740 -280
rect 920 -290 980 -280
rect 1160 -290 1220 -280
rect 1400 -290 1460 -280
rect 1640 -290 1700 -280
rect 1880 -290 1940 -280
rect 2120 -290 2180 -280
rect 2360 -290 2420 -280
rect -130 -350 -40 -290
rect 20 -350 200 -290
rect 260 -350 440 -290
rect 500 -350 680 -290
rect 740 -350 920 -290
rect 980 -350 1160 -290
rect 1220 -350 1400 -290
rect 1460 -350 1640 -290
rect 1700 -350 1880 -290
rect 1940 -350 2120 -290
rect 2180 -350 2360 -290
rect 2420 -350 2680 -290
rect -130 -380 2680 -350
rect 1020 -430 1080 -420
rect 1740 -430 1800 -420
rect -140 -490 1020 -430
rect 1080 -490 1740 -430
rect 1800 -490 2680 -430
rect 1020 -500 1080 -490
rect 1740 -500 1800 -490
rect 1260 -550 1320 -540
rect 1500 -550 1560 -540
rect -140 -610 1260 -550
rect 1320 -610 1500 -550
rect 1560 -610 2680 -550
rect 1260 -620 1320 -610
rect 1500 -620 1560 -610
rect 780 -670 840 -660
rect -140 -730 780 -670
rect 840 -730 2680 -670
rect 780 -740 840 -730
rect 540 -790 600 -780
rect 1980 -790 2040 -780
rect -140 -850 540 -790
rect 600 -850 1980 -790
rect 2040 -850 2680 -790
rect 540 -860 600 -850
rect 1980 -860 2040 -850
rect 60 -910 120 -900
rect 300 -910 360 -900
rect 2220 -910 2280 -900
rect 2460 -910 2520 -900
rect -140 -970 60 -910
rect 120 -970 300 -910
rect 360 -970 2220 -910
rect 2280 -970 2460 -910
rect 2520 -970 2680 -910
rect 60 -980 120 -970
rect 300 -980 360 -970
rect 2220 -980 2280 -970
rect 2460 -980 2520 -970
use sky130_fd_pr__nfet_01v8_lvt_J9Q35V  sky130_fd_pr__nfet_01v8_lvt_J9Q35V_0
array 0 10 -240 0 0 -640
timestamp 1723168442
transform -1 0 88 0 -1 -153
box -88 -107 88 107
use sky130_fd_pr__nfet_01v8_lvt_J9Q35V  sky130_fd_pr__nfet_01v8_lvt_J9Q35V_1
array 0 10 240 0 0 640
timestamp 1723168442
transform 1 0 88 0 1 107
box -88 -107 88 107
<< labels >>
flabel metal2 -140 -610 -80 -550 0 FreeSans 320 0 0 0 D1
port 0 nsew
flabel metal2 -140 -730 -80 -670 0 FreeSans 320 0 0 0 M1
port 1 nsew
flabel metal2 -140 -850 -80 -790 0 FreeSans 320 0 0 0 M2
port 2 nsew
flabel metal2 -140 -970 -80 -910 0 FreeSans 320 0 0 0 M3
port 3 nsew
flabel metal2 -140 -490 -80 -430 0 FreeSans 320 0 0 0 VDDL
port 4 nsew
flabel metal2 -130 -370 -70 -310 0 FreeSans 320 0 0 0 VSS
port 5 nsew
flabel metal2 940 430 1000 490 0 FreeSans 320 0 0 0 MSINK
port 6 nsew
flabel metal1 1170 430 1230 490 0 FreeSans 320 0 0 0 DSINK
port 7 nsew
flabel metal1 1510 420 1570 480 0 FreeSans 320 0 0 0 VG
port 10 nsew
<< end >>
