magic
tech sky130A
magscale 1 2
timestamp 1723401136
<< nwell >>
rect -110 540 550 1120
<< pwell >>
rect -100 -60 550 470
<< metal1 >>
rect -100 1020 500 1120
rect 160 900 240 1020
rect 30 780 400 820
rect 0 680 140 720
rect -40 620 40 680
rect 0 120 40 620
rect 80 500 100 560
rect 160 500 170 560
rect 80 160 120 500
rect 260 380 300 720
rect 360 560 400 780
rect 350 500 360 560
rect 420 500 430 560
rect 230 320 240 380
rect 300 320 310 380
rect 260 300 300 320
rect 200 160 240 260
rect 0 80 200 120
rect 320 40 440 260
rect -100 -60 500 40
<< via1 >>
rect 100 500 160 560
rect 360 500 420 560
rect 240 320 300 380
<< metal2 >>
rect 360 560 420 570
rect 80 500 100 560
rect 160 540 180 560
rect 160 500 360 540
rect 360 490 420 500
rect -100 400 300 440
rect -100 380 -40 400
rect 240 380 300 400
rect 240 310 300 320
use sky130_fd_pr__nfet_01v8_lvt_ZDUAWA  sky130_fd_pr__nfet_01v8_lvt_ZDUAWA_0
timestamp 1723344990
transform 1 0 222 0 1 207
box -275 -260 275 260
use sky130_fd_pr__pfet_01v8_lvt_UT4KY6  sky130_fd_pr__pfet_01v8_lvt_UT4KY6_0
timestamp 1723344990
transform 1 0 192 0 1 831
box -295 -284 295 284
<< labels >>
flabel metal2 -100 380 -40 440 0 FreeSans 800 0 0 0 B
port 1 nsew
flabel metal1 -100 1020 0 1120 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal1 -60 -60 40 40 0 FreeSans 800 0 0 0 VSS
port 4 nsew
flabel metal1 -40 620 20 680 0 FreeSans 800 0 0 0 A
port 0 nsew
flabel metal2 360 500 420 560 0 FreeSans 800 0 0 0 Q
port 2 nsew
<< end >>
