magic
tech sky130A
magscale 1 2
timestamp 1725323004
<< pwell >>
rect -1244 -658 1244 658
<< nnmos >>
rect -1016 -400 -916 400
rect -740 -400 -640 400
rect -464 -400 -364 400
rect -188 -400 -88 400
rect 88 -400 188 400
rect 364 -400 464 400
rect 640 -400 740 400
rect 916 -400 1016 400
<< mvndiff >>
rect -1074 388 -1016 400
rect -1074 -388 -1062 388
rect -1028 -388 -1016 388
rect -1074 -400 -1016 -388
rect -916 388 -858 400
rect -916 -388 -904 388
rect -870 -388 -858 388
rect -916 -400 -858 -388
rect -798 388 -740 400
rect -798 -388 -786 388
rect -752 -388 -740 388
rect -798 -400 -740 -388
rect -640 388 -582 400
rect -640 -388 -628 388
rect -594 -388 -582 388
rect -640 -400 -582 -388
rect -522 388 -464 400
rect -522 -388 -510 388
rect -476 -388 -464 388
rect -522 -400 -464 -388
rect -364 388 -306 400
rect -364 -388 -352 388
rect -318 -388 -306 388
rect -364 -400 -306 -388
rect -246 388 -188 400
rect -246 -388 -234 388
rect -200 -388 -188 388
rect -246 -400 -188 -388
rect -88 388 -30 400
rect -88 -388 -76 388
rect -42 -388 -30 388
rect -88 -400 -30 -388
rect 30 388 88 400
rect 30 -388 42 388
rect 76 -388 88 388
rect 30 -400 88 -388
rect 188 388 246 400
rect 188 -388 200 388
rect 234 -388 246 388
rect 188 -400 246 -388
rect 306 388 364 400
rect 306 -388 318 388
rect 352 -388 364 388
rect 306 -400 364 -388
rect 464 388 522 400
rect 464 -388 476 388
rect 510 -388 522 388
rect 464 -400 522 -388
rect 582 388 640 400
rect 582 -388 594 388
rect 628 -388 640 388
rect 582 -400 640 -388
rect 740 388 798 400
rect 740 -388 752 388
rect 786 -388 798 388
rect 740 -400 798 -388
rect 858 388 916 400
rect 858 -388 870 388
rect 904 -388 916 388
rect 858 -400 916 -388
rect 1016 388 1074 400
rect 1016 -388 1028 388
rect 1062 -388 1074 388
rect 1016 -400 1074 -388
<< mvndiffc >>
rect -1062 -388 -1028 388
rect -904 -388 -870 388
rect -786 -388 -752 388
rect -628 -388 -594 388
rect -510 -388 -476 388
rect -352 -388 -318 388
rect -234 -388 -200 388
rect -76 -388 -42 388
rect 42 -388 76 388
rect 200 -388 234 388
rect 318 -388 352 388
rect 476 -388 510 388
rect 594 -388 628 388
rect 752 -388 786 388
rect 870 -388 904 388
rect 1028 -388 1062 388
<< mvpsubdiff >>
rect -1208 610 1208 622
rect -1208 576 -1100 610
rect 1100 576 1208 610
rect -1208 564 1208 576
rect -1208 514 -1150 564
rect -1208 -514 -1196 514
rect -1162 -514 -1150 514
rect 1150 514 1208 564
rect -1208 -564 -1150 -514
rect 1150 -514 1162 514
rect 1196 -514 1208 514
rect 1150 -564 1208 -514
rect -1208 -576 1208 -564
rect -1208 -610 -1100 -576
rect 1100 -610 1208 -576
rect -1208 -622 1208 -610
<< mvpsubdiffcont >>
rect -1100 576 1100 610
rect -1196 -514 -1162 514
rect 1162 -514 1196 514
rect -1100 -610 1100 -576
<< poly >>
rect -1016 472 -916 488
rect -1016 438 -1000 472
rect -932 438 -916 472
rect -1016 400 -916 438
rect -740 472 -640 488
rect -740 438 -724 472
rect -656 438 -640 472
rect -740 400 -640 438
rect -464 472 -364 488
rect -464 438 -448 472
rect -380 438 -364 472
rect -464 400 -364 438
rect -188 472 -88 488
rect -188 438 -172 472
rect -104 438 -88 472
rect -188 400 -88 438
rect 88 472 188 488
rect 88 438 104 472
rect 172 438 188 472
rect 88 400 188 438
rect 364 472 464 488
rect 364 438 380 472
rect 448 438 464 472
rect 364 400 464 438
rect 640 472 740 488
rect 640 438 656 472
rect 724 438 740 472
rect 640 400 740 438
rect 916 472 1016 488
rect 916 438 932 472
rect 1000 438 1016 472
rect 916 400 1016 438
rect -1016 -438 -916 -400
rect -1016 -472 -1000 -438
rect -932 -472 -916 -438
rect -1016 -488 -916 -472
rect -740 -438 -640 -400
rect -740 -472 -724 -438
rect -656 -472 -640 -438
rect -740 -488 -640 -472
rect -464 -438 -364 -400
rect -464 -472 -448 -438
rect -380 -472 -364 -438
rect -464 -488 -364 -472
rect -188 -438 -88 -400
rect -188 -472 -172 -438
rect -104 -472 -88 -438
rect -188 -488 -88 -472
rect 88 -438 188 -400
rect 88 -472 104 -438
rect 172 -472 188 -438
rect 88 -488 188 -472
rect 364 -438 464 -400
rect 364 -472 380 -438
rect 448 -472 464 -438
rect 364 -488 464 -472
rect 640 -438 740 -400
rect 640 -472 656 -438
rect 724 -472 740 -438
rect 640 -488 740 -472
rect 916 -438 1016 -400
rect 916 -472 932 -438
rect 1000 -472 1016 -438
rect 916 -488 1016 -472
<< polycont >>
rect -1000 438 -932 472
rect -724 438 -656 472
rect -448 438 -380 472
rect -172 438 -104 472
rect 104 438 172 472
rect 380 438 448 472
rect 656 438 724 472
rect 932 438 1000 472
rect -1000 -472 -932 -438
rect -724 -472 -656 -438
rect -448 -472 -380 -438
rect -172 -472 -104 -438
rect 104 -472 172 -438
rect 380 -472 448 -438
rect 656 -472 724 -438
rect 932 -472 1000 -438
<< locali >>
rect -1196 576 -1100 610
rect 1100 576 1196 610
rect -1196 514 -1162 576
rect 1162 514 1196 576
rect -1016 438 -1000 472
rect -932 438 -916 472
rect -740 438 -724 472
rect -656 438 -640 472
rect -464 438 -448 472
rect -380 438 -364 472
rect -188 438 -172 472
rect -104 438 -88 472
rect 88 438 104 472
rect 172 438 188 472
rect 364 438 380 472
rect 448 438 464 472
rect 640 438 656 472
rect 724 438 740 472
rect 916 438 932 472
rect 1000 438 1016 472
rect -1062 388 -1028 404
rect -1062 -404 -1028 -388
rect -904 388 -870 404
rect -904 -404 -870 -388
rect -786 388 -752 404
rect -786 -404 -752 -388
rect -628 388 -594 404
rect -628 -404 -594 -388
rect -510 388 -476 404
rect -510 -404 -476 -388
rect -352 388 -318 404
rect -352 -404 -318 -388
rect -234 388 -200 404
rect -234 -404 -200 -388
rect -76 388 -42 404
rect -76 -404 -42 -388
rect 42 388 76 404
rect 42 -404 76 -388
rect 200 388 234 404
rect 200 -404 234 -388
rect 318 388 352 404
rect 318 -404 352 -388
rect 476 388 510 404
rect 476 -404 510 -388
rect 594 388 628 404
rect 594 -404 628 -388
rect 752 388 786 404
rect 752 -404 786 -388
rect 870 388 904 404
rect 870 -404 904 -388
rect 1028 388 1062 404
rect 1028 -404 1062 -388
rect -1016 -472 -1000 -438
rect -932 -472 -916 -438
rect -740 -472 -724 -438
rect -656 -472 -640 -438
rect -464 -472 -448 -438
rect -380 -472 -364 -438
rect -188 -472 -172 -438
rect -104 -472 -88 -438
rect 88 -472 104 -438
rect 172 -472 188 -438
rect 364 -472 380 -438
rect 448 -472 464 -438
rect 640 -472 656 -438
rect 724 -472 740 -438
rect 916 -472 932 -438
rect 1000 -472 1016 -438
rect -1196 -576 -1162 -514
rect 1162 -576 1196 -514
rect -1196 -610 -1100 -576
rect 1100 -610 1196 -576
<< viali >>
rect -1000 438 -932 472
rect -724 438 -656 472
rect -448 438 -380 472
rect -172 438 -104 472
rect 104 438 172 472
rect 380 438 448 472
rect 656 438 724 472
rect 932 438 1000 472
rect -1196 -230 -1162 230
rect -1062 -371 -1028 -61
rect -904 61 -870 371
rect -786 61 -752 371
rect -628 -371 -594 -61
rect -510 -371 -476 -61
rect -352 61 -318 371
rect -234 61 -200 371
rect -76 -371 -42 -61
rect 42 -371 76 -61
rect 200 61 234 371
rect 318 61 352 371
rect 476 -371 510 -61
rect 594 -371 628 -61
rect 752 61 786 371
rect 870 61 904 371
rect 1028 -371 1062 -61
rect 1162 -230 1196 230
rect -1000 -472 -932 -438
rect -724 -472 -656 -438
rect -448 -472 -380 -438
rect -172 -472 -104 -438
rect 104 -472 172 -438
rect 380 -472 448 -438
rect 656 -472 724 -438
rect 932 -472 1000 -438
rect -465 -610 465 -576
<< metal1 >>
rect -1012 472 -920 478
rect -1012 438 -1000 472
rect -932 438 -920 472
rect -1012 432 -920 438
rect -736 472 -644 478
rect -736 438 -724 472
rect -656 438 -644 472
rect -736 432 -644 438
rect -460 472 -368 478
rect -460 438 -448 472
rect -380 438 -368 472
rect -460 432 -368 438
rect -184 472 -92 478
rect -184 438 -172 472
rect -104 438 -92 472
rect -184 432 -92 438
rect 92 472 184 478
rect 92 438 104 472
rect 172 438 184 472
rect 92 432 184 438
rect 368 472 460 478
rect 368 438 380 472
rect 448 438 460 472
rect 368 432 460 438
rect 644 472 736 478
rect 644 438 656 472
rect 724 438 736 472
rect 644 432 736 438
rect 920 472 1012 478
rect 920 438 932 472
rect 1000 438 1012 472
rect 920 432 1012 438
rect -910 371 -864 383
rect -1202 230 -1156 242
rect -1202 -230 -1196 230
rect -1162 -230 -1156 230
rect -910 61 -904 371
rect -870 61 -864 371
rect -910 49 -864 61
rect -792 371 -746 383
rect -792 61 -786 371
rect -752 61 -746 371
rect -792 49 -746 61
rect -358 371 -312 383
rect -358 61 -352 371
rect -318 61 -312 371
rect -358 49 -312 61
rect -240 371 -194 383
rect -240 61 -234 371
rect -200 61 -194 371
rect -240 49 -194 61
rect 194 371 240 383
rect 194 61 200 371
rect 234 61 240 371
rect 194 49 240 61
rect 312 371 358 383
rect 312 61 318 371
rect 352 61 358 371
rect 312 49 358 61
rect 746 371 792 383
rect 746 61 752 371
rect 786 61 792 371
rect 746 49 792 61
rect 864 371 910 383
rect 864 61 870 371
rect 904 61 910 371
rect 864 49 910 61
rect 1156 230 1202 242
rect -1202 -242 -1156 -230
rect -1068 -61 -1022 -49
rect -1068 -371 -1062 -61
rect -1028 -371 -1022 -61
rect -1068 -383 -1022 -371
rect -634 -61 -588 -49
rect -634 -371 -628 -61
rect -594 -371 -588 -61
rect -634 -383 -588 -371
rect -516 -61 -470 -49
rect -516 -371 -510 -61
rect -476 -371 -470 -61
rect -516 -383 -470 -371
rect -82 -61 -36 -49
rect -82 -371 -76 -61
rect -42 -371 -36 -61
rect -82 -383 -36 -371
rect 36 -61 82 -49
rect 36 -371 42 -61
rect 76 -371 82 -61
rect 36 -383 82 -371
rect 470 -61 516 -49
rect 470 -371 476 -61
rect 510 -371 516 -61
rect 470 -383 516 -371
rect 588 -61 634 -49
rect 588 -371 594 -61
rect 628 -371 634 -61
rect 588 -383 634 -371
rect 1022 -61 1068 -49
rect 1022 -371 1028 -61
rect 1062 -371 1068 -61
rect 1156 -230 1162 230
rect 1196 -230 1202 230
rect 1156 -242 1202 -230
rect 1022 -383 1068 -371
rect -1012 -438 -920 -432
rect -1012 -472 -1000 -438
rect -932 -472 -920 -438
rect -1012 -478 -920 -472
rect -736 -438 -644 -432
rect -736 -472 -724 -438
rect -656 -472 -644 -438
rect -736 -478 -644 -472
rect -460 -438 -368 -432
rect -460 -472 -448 -438
rect -380 -472 -368 -438
rect -460 -478 -368 -472
rect -184 -438 -92 -432
rect -184 -472 -172 -438
rect -104 -472 -92 -438
rect -184 -478 -92 -472
rect 92 -438 184 -432
rect 92 -472 104 -438
rect 172 -472 184 -438
rect 92 -478 184 -472
rect 368 -438 460 -432
rect 368 -472 380 -438
rect 448 -472 460 -438
rect 368 -478 460 -472
rect 644 -438 736 -432
rect 644 -472 656 -438
rect 724 -472 736 -438
rect 644 -478 736 -472
rect 920 -438 1012 -432
rect 920 -472 932 -438
rect 1000 -472 1012 -438
rect 920 -478 1012 -472
rect -477 -576 477 -570
rect -477 -610 -465 -576
rect 465 -610 477 -576
rect -477 -616 477 -610
<< properties >>
string FIXED_BBOX -1179 -593 1179 593
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 4 l 0.50 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 40 viagr 40 viagl 40 viagt 0
string sky130_fd_pr__nfet_03v3_nvt_7WRH84 parameters
<< end >>
