magic
tech sky130A
magscale 1 2
timestamp 1713067979
<< locali >>
rect 1640 1620 5180 1780
rect 1520 880 5320 900
rect 1520 780 5340 880
rect 1520 760 5320 780
rect 1520 700 4080 760
rect 1520 -1120 1660 700
rect 2920 -280 4060 700
rect 2920 -920 3120 -280
rect 3860 -920 4060 -280
rect 2920 -1120 4060 -920
rect 1520 -1260 5320 -1120
<< metal1 >>
rect 1640 1620 5180 1780
rect 2180 1440 2280 1620
rect 2700 1440 2800 1620
rect 3980 1440 4080 1620
rect 4480 1440 4580 1620
rect 1640 1220 3080 1400
rect 3740 1220 5180 1400
rect 1780 1060 4940 1180
rect 1520 880 1660 900
rect 1520 760 5300 880
rect 1520 700 4080 760
rect 1520 -1120 1660 700
rect 3840 -140 4060 -120
rect 2900 -280 4060 -140
rect 1960 -440 2080 -420
rect 1960 -700 2000 -440
rect 2060 -700 2080 -440
rect 1960 -720 2080 -700
rect 2480 -440 2600 -420
rect 2480 -700 2500 -440
rect 2560 -700 2600 -440
rect 2480 -720 2600 -700
rect 2900 -1120 3120 -280
rect 3180 -440 3280 -420
rect 3180 -700 3200 -440
rect 3260 -700 3280 -440
rect 3440 -700 3540 -280
rect 3700 -440 3800 -420
rect 3760 -700 3800 -440
rect 3180 -720 3280 -700
rect 3700 -720 3800 -700
rect 3840 -1120 4060 -280
rect 4380 -440 4480 -420
rect 4440 -700 4480 -440
rect 4380 -720 4480 -700
rect 4900 -440 5000 -420
rect 4960 -700 5000 -440
rect 4900 -720 5000 -700
rect 1520 -1260 5320 -1120
<< via1 >>
rect 2000 -700 2060 -440
rect 2500 -700 2560 -440
rect 3200 -700 3260 -440
rect 3700 -700 3760 -440
rect 4380 -700 4440 -440
rect 4900 -700 4960 -440
<< metal2 >>
rect 1960 -440 5020 -420
rect 1960 -700 2000 -440
rect 2060 -700 2500 -440
rect 2560 -700 3200 -440
rect 3260 -700 3700 -440
rect 3760 -700 4380 -440
rect 4440 -700 4900 -440
rect 4960 -700 5020 -440
rect 1960 -720 5020 -700
use sky130_fd_pr__nfet_01v8_5WCAAQ  sky130_fd_pr__nfet_01v8_5WCAAQ_0
timestamp 1713067979
transform -1 0 2283 0 1 -221
box -683 -979 683 979
use sky130_fd_pr__nfet_01v8_33LZYU  sky130_fd_pr__nfet_01v8_33LZYU_0
timestamp 1713067979
transform 1 0 3485 0 1 -581
box -425 -379 425 379
use sky130_fd_pr__nfet_01v8_MM2THM  sky130_fd_pr__nfet_01v8_MM2THM_0
timestamp 1713067979
transform 1 0 4683 0 1 -190
box -683 -1010 683 1010
use sky130_fd_pr__pfet_01v8_D6KM8H  sky130_fd_pr__pfet_01v8_D6KM8H_0
timestamp 1713067979
transform 1 0 2483 0 1 1384
box -683 -384 683 384
use sky130_fd_pr__pfet_01v8_D6KM8H  sky130_fd_pr__pfet_01v8_D6KM8H_1
timestamp 1713067979
transform 1 0 4283 0 1 1384
box -683 -384 683 384
<< end >>
