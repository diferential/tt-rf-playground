magic
tech sky130A
timestamp 1720664591
<< metal2 >>
rect 0 -135 20 155
rect 85 135 145 155
rect 535 135 595 155
rect 985 135 1045 155
rect 1435 -115 1455 155
rect 305 -135 365 -115
rect 755 -135 815 -115
rect 1195 -135 1255 -115
rect 1340 -135 1455 -115
use pll_inv1  pll_inv1_0
array 0 2 -450 0 0 -290
timestamp 1720664591
transform -1 0 400 0 -1 -25
box -50 -45 400 245
use pll_inv1  pll_inv1_1
array 0 3 450 0 0 290
timestamp 1720664591
transform 1 0 50 0 1 45
box -50 -45 400 245
<< end >>
