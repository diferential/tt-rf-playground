magic
tech sky130A
magscale 1 2
timestamp 1719784689
<< error_p >>
rect 191 -286 249 -280
rect 191 -320 203 -286
rect 191 -326 249 -320
rect 200 -460 205 -450
rect 235 -460 240 -450
<< error_s >>
rect 3724 870 3732 970
rect 3752 890 3760 970
rect 3724 610 3732 710
rect 3752 630 3760 710
rect 3724 350 3732 450
rect 3752 370 3760 450
rect 5709 -407 5767 -401
rect 5709 -441 5721 -407
rect 5709 -447 5767 -441
rect 5563 -690 5574 -546
rect 5709 -601 5767 -595
rect 5709 -635 5721 -601
rect 5709 -641 5767 -635
<< pwell >>
rect -11640 -11730 20630 9310
<< nmos >>
rect 4780 210 4810 300
rect 4890 210 4920 300
rect 5000 210 5030 300
rect 4780 -80 4810 10
rect 4890 -80 4920 10
rect 5000 -80 5030 10
rect 5390 -200 5420 0
rect 480 -300 520 -200
rect 620 -300 660 -200
rect 760 -300 800 -200
rect 900 -300 940 -200
rect 1040 -300 1080 -200
rect 1180 -300 1220 -200
rect 205 -442 235 -358
rect 480 -460 520 -360
rect 620 -460 660 -360
rect 760 -460 800 -360
rect 900 -460 940 -360
rect 1040 -460 1080 -360
rect 1180 -460 1220 -360
rect 4670 -690 4700 -600
rect 4780 -690 4810 -600
rect 4860 -690 4890 -600
rect 4970 -690 5000 -600
rect 5050 -690 5080 -600
rect 5160 -690 5190 -600
rect 1430 -1550 1470 -1460
rect 1520 -1550 1560 -1460
rect 1610 -1550 1650 -1460
rect 1700 -1550 1740 -1460
rect 1900 -1550 1940 -1460
rect 1990 -1550 2030 -1460
rect 2080 -1550 2120 -1460
rect 2170 -1550 2210 -1460
rect 2370 -1550 2410 -1460
rect 2460 -1550 2500 -1460
rect 2550 -1550 2590 -1460
rect 2640 -1550 2680 -1460
rect 1430 -1700 1470 -1610
rect 1520 -1700 1560 -1610
rect 1610 -1700 1650 -1610
rect 1700 -1700 1740 -1610
rect 1900 -1700 1940 -1610
rect 1990 -1700 2030 -1610
rect 2080 -1700 2120 -1610
rect 2170 -1700 2210 -1610
rect 2370 -1700 2410 -1610
rect 2460 -1700 2500 -1610
rect 2550 -1700 2590 -1610
rect 2640 -1700 2680 -1610
rect 3720 -1710 3750 -1620
rect 1430 -1850 1470 -1760
rect 1520 -1850 1560 -1760
rect 1610 -1850 1650 -1760
rect 1700 -1850 1740 -1760
rect 1900 -1850 1940 -1760
rect 1990 -1850 2030 -1760
rect 2080 -1850 2120 -1760
rect 2170 -1850 2210 -1760
rect 2370 -1850 2410 -1760
rect 2460 -1850 2500 -1760
rect 2550 -1850 2590 -1760
rect 2640 -1850 2680 -1760
rect 3640 -1910 3670 -1820
rect 3720 -1910 3750 -1820
rect 4030 -1910 4060 -1820
rect 4140 -1910 4170 -1820
rect 4220 -1910 4250 -1820
rect 1430 -2000 1470 -1910
rect 1520 -2000 1560 -1910
rect 1610 -2000 1650 -1910
rect 1700 -2000 1740 -1910
rect 1900 -2000 1940 -1910
rect 1990 -2000 2030 -1910
rect 2080 -2000 2120 -1910
rect 2170 -2000 2210 -1910
rect 2370 -2000 2410 -1910
rect 2460 -2000 2500 -1910
rect 2550 -2000 2590 -1910
rect 2640 -2000 2680 -1910
rect 1430 -2150 1470 -2060
rect 1520 -2150 1560 -2060
rect 1610 -2150 1650 -2060
rect 1700 -2150 1740 -2060
rect 1900 -2150 1940 -2060
rect 1990 -2150 2030 -2060
rect 2080 -2150 2120 -2060
rect 2170 -2150 2210 -2060
rect 2370 -2150 2410 -2060
rect 2460 -2150 2500 -2060
rect 2550 -2150 2590 -2060
rect 2640 -2150 2680 -2060
rect 1430 -2300 1470 -2210
rect 1520 -2300 1560 -2210
rect 1610 -2300 1650 -2210
rect 1700 -2300 1740 -2210
rect 1900 -2300 1940 -2210
rect 1990 -2300 2030 -2210
rect 2080 -2300 2120 -2210
rect 2170 -2300 2210 -2210
rect 2370 -2300 2410 -2210
rect 2460 -2300 2500 -2210
rect 2550 -2300 2590 -2210
rect 2640 -2300 2680 -2210
<< ndiff >>
rect 4710 280 4780 300
rect 4710 230 4720 280
rect 4760 230 4780 280
rect 4710 210 4780 230
rect 4810 270 4890 300
rect 4810 230 4830 270
rect 4870 230 4890 270
rect 4810 210 4890 230
rect 4920 210 5000 300
rect 5030 280 5100 300
rect 5030 240 5050 280
rect 5090 240 5100 280
rect 5030 210 5100 240
rect 4710 -20 4780 10
rect 4710 -60 4720 -20
rect 4760 -60 4780 -20
rect 4710 -80 4780 -60
rect 4810 -80 4890 10
rect 4920 -20 5000 10
rect 4920 -60 4940 -20
rect 4980 -60 5000 -20
rect 4920 -80 5000 -60
rect 5030 -20 5100 10
rect 5030 -60 5050 -20
rect 5090 -60 5100 -20
rect 5030 -80 5100 -60
rect 5320 -80 5390 0
rect 5320 -120 5330 -80
rect 5370 -120 5390 -80
rect 5320 -200 5390 -120
rect 5420 -200 5470 0
rect 380 -220 480 -200
rect 380 -280 400 -220
rect 460 -280 480 -220
rect 380 -300 480 -280
rect 520 -220 620 -200
rect 520 -280 540 -220
rect 600 -280 620 -220
rect 520 -300 620 -280
rect 660 -220 760 -200
rect 660 -280 680 -220
rect 740 -280 760 -220
rect 660 -300 760 -280
rect 800 -220 900 -200
rect 800 -280 820 -220
rect 880 -280 900 -220
rect 800 -300 900 -280
rect 940 -220 1040 -200
rect 940 -280 960 -220
rect 1020 -280 1040 -220
rect 940 -300 1040 -280
rect 1080 -220 1180 -200
rect 1080 -280 1100 -220
rect 1160 -280 1180 -220
rect 1080 -300 1180 -280
rect 1220 -220 1320 -200
rect 1220 -280 1240 -220
rect 1300 -280 1320 -220
rect 1220 -300 1320 -280
rect 147 -360 205 -358
rect 140 -370 205 -360
rect 140 -430 159 -370
rect 193 -430 205 -370
rect 140 -440 205 -430
rect 147 -442 205 -440
rect 235 -370 293 -358
rect 235 -430 247 -370
rect 281 -430 293 -370
rect 235 -442 293 -430
rect 380 -380 480 -360
rect 380 -440 400 -380
rect 460 -440 480 -380
rect 380 -460 480 -440
rect 520 -380 620 -360
rect 520 -440 540 -380
rect 600 -440 620 -380
rect 520 -460 620 -440
rect 660 -380 760 -360
rect 660 -440 680 -380
rect 740 -440 760 -380
rect 660 -460 760 -440
rect 800 -380 900 -360
rect 800 -440 820 -380
rect 880 -440 900 -380
rect 800 -460 900 -440
rect 940 -380 1040 -360
rect 940 -440 960 -380
rect 1020 -440 1040 -380
rect 940 -460 1040 -440
rect 1080 -380 1180 -360
rect 1080 -440 1100 -380
rect 1160 -440 1180 -380
rect 1080 -460 1180 -440
rect 1220 -380 1320 -360
rect 1220 -440 1240 -380
rect 1300 -440 1320 -380
rect 1220 -460 1320 -440
rect 4600 -620 4670 -600
rect 4600 -660 4610 -620
rect 4650 -660 4670 -620
rect 4600 -690 4670 -660
rect 4700 -620 4780 -600
rect 4700 -660 4720 -620
rect 4760 -660 4780 -620
rect 4700 -690 4780 -660
rect 4810 -690 4860 -600
rect 4890 -620 4970 -600
rect 4890 -660 4910 -620
rect 4950 -660 4970 -620
rect 4890 -690 4970 -660
rect 5000 -690 5050 -600
rect 5080 -630 5160 -600
rect 5080 -670 5100 -630
rect 5140 -670 5160 -630
rect 5080 -690 5160 -670
rect 5190 -630 5260 -600
rect 5190 -670 5210 -630
rect 5250 -670 5260 -630
rect 5190 -690 5260 -670
rect 5320 -690 5520 -600
rect 1380 -1550 1430 -1460
rect 1470 -1550 1520 -1460
rect 1560 -1550 1610 -1460
rect 1650 -1550 1700 -1460
rect 1740 -1550 1790 -1460
rect 1850 -1550 1900 -1460
rect 1940 -1550 1990 -1460
rect 2030 -1550 2080 -1460
rect 2120 -1550 2170 -1460
rect 2210 -1550 2260 -1460
rect 2320 -1550 2370 -1460
rect 2410 -1550 2460 -1460
rect 2500 -1550 2550 -1460
rect 2590 -1550 2640 -1460
rect 2680 -1550 2730 -1460
rect 1380 -1700 1430 -1610
rect 1470 -1700 1520 -1610
rect 1560 -1700 1610 -1610
rect 1650 -1700 1700 -1610
rect 1740 -1700 1790 -1610
rect 1850 -1700 1900 -1610
rect 1940 -1700 1990 -1610
rect 2030 -1700 2080 -1610
rect 2120 -1700 2170 -1610
rect 2210 -1700 2260 -1610
rect 2320 -1700 2370 -1610
rect 2410 -1700 2460 -1610
rect 2500 -1700 2550 -1610
rect 2590 -1700 2640 -1610
rect 2680 -1700 2730 -1610
rect 3770 -1620 3810 -1550
rect 3650 -1710 3720 -1620
rect 3750 -1710 3810 -1620
rect 1380 -1850 1430 -1760
rect 1470 -1850 1520 -1760
rect 1560 -1850 1610 -1760
rect 1650 -1850 1700 -1760
rect 1740 -1850 1790 -1760
rect 1850 -1850 1900 -1760
rect 1940 -1850 1990 -1760
rect 2030 -1850 2080 -1760
rect 2120 -1850 2170 -1760
rect 2210 -1850 2260 -1760
rect 2320 -1850 2370 -1760
rect 2410 -1850 2460 -1760
rect 2500 -1850 2550 -1760
rect 2590 -1850 2640 -1760
rect 2680 -1850 2730 -1760
rect 3770 -1820 3810 -1710
rect 4080 -1820 4120 -1730
rect 3570 -1910 3640 -1820
rect 3670 -1910 3720 -1820
rect 3750 -1910 3810 -1820
rect 3960 -1910 4030 -1820
rect 4060 -1910 4140 -1820
rect 4170 -1910 4220 -1820
rect 4250 -1910 4320 -1820
rect 1380 -2000 1430 -1910
rect 1470 -2000 1520 -1910
rect 1560 -2000 1610 -1910
rect 1650 -2000 1700 -1910
rect 1740 -2000 1790 -1910
rect 1850 -2000 1900 -1910
rect 1940 -2000 1990 -1910
rect 2030 -2000 2080 -1910
rect 2120 -2000 2170 -1910
rect 2210 -2000 2260 -1910
rect 2320 -2000 2370 -1910
rect 2410 -2000 2460 -1910
rect 2500 -2000 2550 -1910
rect 2590 -2000 2640 -1910
rect 2680 -2000 2730 -1910
rect 3770 -1970 3810 -1910
rect 4080 -1940 4120 -1910
rect 1380 -2150 1430 -2060
rect 1470 -2150 1520 -2060
rect 1560 -2150 1610 -2060
rect 1650 -2150 1700 -2060
rect 1740 -2150 1790 -2060
rect 1850 -2150 1900 -2060
rect 1940 -2150 1990 -2060
rect 2030 -2150 2080 -2060
rect 2120 -2150 2170 -2060
rect 2210 -2150 2260 -2060
rect 2320 -2150 2370 -2060
rect 2410 -2150 2460 -2060
rect 2500 -2150 2550 -2060
rect 2590 -2150 2640 -2060
rect 2680 -2150 2730 -2060
rect 1380 -2300 1430 -2210
rect 1470 -2300 1520 -2210
rect 1560 -2300 1610 -2210
rect 1650 -2300 1700 -2210
rect 1740 -2300 1790 -2210
rect 1850 -2300 1900 -2210
rect 1940 -2300 1990 -2210
rect 2030 -2300 2080 -2210
rect 2120 -2300 2170 -2210
rect 2210 -2300 2260 -2210
rect 2320 -2300 2370 -2210
rect 2410 -2300 2460 -2210
rect 2500 -2300 2550 -2210
rect 2590 -2300 2640 -2210
rect 2680 -2300 2730 -2210
<< ndiffc >>
rect 4720 230 4760 280
rect 4830 230 4870 270
rect 5050 240 5090 280
rect 4720 -60 4760 -20
rect 4940 -60 4980 -20
rect 5050 -60 5090 -20
rect 5330 -120 5370 -80
rect 400 -280 460 -220
rect 540 -280 600 -220
rect 680 -280 740 -220
rect 820 -280 880 -220
rect 960 -280 1020 -220
rect 1100 -280 1160 -220
rect 1240 -280 1300 -220
rect 159 -430 193 -370
rect 247 -430 281 -370
rect 400 -440 460 -380
rect 540 -440 600 -380
rect 680 -440 740 -380
rect 820 -440 880 -380
rect 960 -440 1020 -380
rect 1100 -440 1160 -380
rect 1240 -440 1300 -380
rect 4610 -660 4650 -620
rect 4720 -660 4760 -620
rect 4910 -660 4950 -620
rect 5100 -670 5140 -630
rect 5210 -670 5250 -630
<< poly >>
rect 4780 300 4810 330
rect 4890 300 4920 330
rect 5000 300 5030 330
rect 4780 180 4810 210
rect 4890 180 4920 210
rect 5000 190 5030 210
rect 4970 160 5100 190
rect 4710 100 4840 130
rect 4710 60 4720 100
rect 4760 60 4840 100
rect 4970 120 5050 160
rect 5090 120 5100 160
rect 4970 90 5100 120
rect 4710 30 4840 60
rect 4780 10 4810 30
rect 4890 10 4920 40
rect 5000 10 5030 40
rect 200 -80 1800 -40
rect 5390 0 5420 30
rect 4780 -110 4810 -80
rect 4890 -110 4920 -80
rect 5000 -110 5030 -80
rect 480 -200 520 -160
rect 620 -200 660 -160
rect 760 -200 800 -160
rect 900 -200 940 -160
rect 1040 -200 1080 -160
rect 1180 -200 1220 -160
rect 187 -286 253 -270
rect 187 -320 203 -286
rect 237 -320 253 -286
rect 5390 -230 5420 -200
rect 187 -336 253 -320
rect 205 -358 235 -336
rect 40 -460 120 -360
rect 480 -360 520 -300
rect 620 -360 660 -300
rect 760 -360 800 -300
rect 900 -360 940 -300
rect 1040 -360 1080 -300
rect 1180 -360 1220 -300
rect 205 -460 235 -442
rect 200 -480 240 -460
rect 480 -520 520 -460
rect 620 -520 660 -460
rect 760 -520 800 -460
rect 900 -520 940 -460
rect 1040 -520 1080 -460
rect 1180 -520 1220 -460
rect 4670 -600 4700 -450
rect 4780 -600 4810 -450
rect 4940 -510 5000 -490
rect 4940 -550 4950 -510
rect 4990 -550 5000 -510
rect 4940 -570 5000 -550
rect 4860 -600 4890 -570
rect 4970 -600 5000 -570
rect 5050 -600 5080 -450
rect 5160 -600 5190 -450
rect 520 -720 620 -620
rect 4670 -790 4700 -690
rect 4780 -790 4810 -690
rect 4860 -710 4890 -690
rect 4860 -730 4920 -710
rect 4970 -720 5000 -690
rect 4860 -770 4870 -730
rect 4910 -770 4920 -730
rect 4860 -790 4920 -770
rect 5050 -790 5080 -690
rect 5160 -790 5190 -690
rect 1430 -1460 1470 -1400
rect 1520 -1460 1560 -1400
rect 1610 -1460 1650 -1400
rect 1700 -1460 1740 -1400
rect 1900 -1460 1940 -1400
rect 1990 -1460 2030 -1400
rect 2080 -1460 2120 -1400
rect 2170 -1460 2210 -1400
rect 2370 -1460 2410 -1400
rect 2460 -1460 2500 -1400
rect 2550 -1460 2590 -1400
rect 2640 -1460 2680 -1400
rect 1430 -1610 1470 -1550
rect 1520 -1610 1560 -1550
rect 1610 -1610 1650 -1550
rect 1700 -1610 1740 -1550
rect 1900 -1610 1940 -1550
rect 1990 -1610 2030 -1550
rect 2080 -1610 2120 -1550
rect 2170 -1610 2210 -1550
rect 2370 -1610 2410 -1550
rect 2460 -1610 2500 -1550
rect 2550 -1610 2590 -1550
rect 2640 -1610 2680 -1550
rect 1430 -1760 1470 -1700
rect 1520 -1760 1560 -1700
rect 1610 -1760 1650 -1700
rect 1700 -1760 1740 -1700
rect 1900 -1760 1940 -1700
rect 1990 -1760 2030 -1700
rect 2080 -1760 2120 -1700
rect 2170 -1760 2210 -1700
rect 2370 -1760 2410 -1700
rect 2460 -1760 2500 -1700
rect 2550 -1760 2590 -1700
rect 2640 -1760 2680 -1700
rect 3570 -1730 3630 -1600
rect 3720 -1620 3750 -1590
rect 3570 -1800 3670 -1730
rect 3720 -1740 3750 -1710
rect 3640 -1820 3670 -1800
rect 3720 -1820 3750 -1790
rect 4030 -1820 4060 -1790
rect 4140 -1820 4170 -1790
rect 4220 -1800 4370 -1770
rect 4220 -1820 4250 -1800
rect 1430 -1910 1470 -1850
rect 1520 -1910 1560 -1850
rect 1610 -1910 1650 -1850
rect 1700 -1910 1740 -1850
rect 1900 -1910 1940 -1850
rect 1990 -1910 2030 -1850
rect 2080 -1910 2120 -1850
rect 2170 -1910 2210 -1850
rect 2370 -1910 2410 -1850
rect 2460 -1910 2500 -1850
rect 2550 -1910 2590 -1850
rect 2640 -1910 2680 -1850
rect 3640 -1940 3670 -1910
rect 3720 -1940 3750 -1910
rect 4030 -1940 4060 -1910
rect 4140 -1940 4170 -1910
rect 4220 -1940 4250 -1910
rect 4340 -1940 4370 -1800
rect 1430 -2060 1470 -2000
rect 1520 -2060 1560 -2000
rect 1610 -2060 1650 -2000
rect 1700 -2060 1740 -2000
rect 1900 -2060 1940 -2000
rect 1990 -2060 2030 -2000
rect 2080 -2060 2120 -2000
rect 2170 -2060 2210 -2000
rect 2370 -2060 2410 -2000
rect 2460 -2060 2500 -2000
rect 2550 -2060 2590 -2000
rect 2640 -2060 2680 -2000
rect 1430 -2210 1470 -2150
rect 1520 -2210 1560 -2150
rect 1610 -2210 1650 -2150
rect 1700 -2210 1740 -2150
rect 1900 -2210 1940 -2150
rect 1990 -2210 2030 -2150
rect 2080 -2210 2120 -2150
rect 2170 -2210 2210 -2150
rect 2370 -2210 2410 -2150
rect 2460 -2210 2500 -2150
rect 2550 -2210 2590 -2150
rect 2640 -2210 2680 -2150
rect 1430 -2360 1470 -2300
rect 1520 -2360 1560 -2300
rect 1610 -2360 1650 -2300
rect 1700 -2360 1740 -2300
rect 1900 -2360 1940 -2300
rect 1990 -2360 2030 -2300
rect 2080 -2360 2120 -2300
rect 2170 -2360 2210 -2300
rect 2370 -2360 2410 -2300
rect 2460 -2360 2500 -2300
rect 2550 -2360 2590 -2300
rect 2640 -2360 2680 -2300
<< polycont >>
rect 4720 60 4760 100
rect 5050 120 5090 160
rect 203 -320 237 -286
rect 4950 -550 4990 -510
rect 4870 -770 4910 -730
<< locali >>
rect 4720 280 4760 300
rect 4720 210 4760 230
rect 4830 270 4870 300
rect 4830 210 4870 230
rect 5050 280 5090 300
rect 5050 220 5090 240
rect 5050 160 5090 180
rect 4720 100 4760 130
rect 5050 100 5090 120
rect 4720 40 4760 60
rect 4720 -20 4760 0
rect 200 -80 1800 -40
rect 4720 -80 4760 -60
rect 4940 -20 4980 10
rect 4940 -80 4980 -60
rect 5050 -20 5090 10
rect 5330 -20 5390 20
rect 5050 -80 5090 -60
rect 5330 -80 5370 -60
rect 5330 -140 5370 -120
rect 5510 -80 5710 0
rect 5510 -120 5590 -80
rect 5630 -120 5710 -80
rect 5510 -200 5710 -120
rect 5770 -80 5810 -60
rect 5770 -140 5810 -120
rect 380 -220 480 -200
rect 380 -280 400 -220
rect 460 -280 480 -220
rect 187 -320 203 -286
rect 237 -320 253 -286
rect 380 -300 480 -280
rect 520 -220 620 -200
rect 520 -280 540 -220
rect 600 -280 620 -220
rect 520 -300 620 -280
rect 660 -220 760 -200
rect 660 -280 680 -220
rect 740 -280 760 -220
rect 660 -300 760 -280
rect 800 -220 900 -200
rect 800 -280 820 -220
rect 880 -280 900 -220
rect 800 -300 900 -280
rect 940 -220 1040 -200
rect 940 -280 960 -220
rect 1020 -280 1040 -220
rect 940 -300 1040 -280
rect 1080 -220 1180 -200
rect 1080 -280 1100 -220
rect 1160 -280 1180 -220
rect 1080 -300 1180 -280
rect 1220 -220 1320 -200
rect 1220 -280 1240 -220
rect 1300 -280 1320 -220
rect 1220 -300 1320 -280
rect 159 -360 193 -354
rect 40 -370 193 -360
rect 40 -380 159 -370
rect 40 -440 60 -380
rect 120 -430 159 -380
rect 120 -440 193 -430
rect 40 -460 120 -440
rect 159 -446 193 -440
rect 247 -370 281 -354
rect 247 -446 281 -430
rect 380 -380 480 -350
rect 380 -440 400 -380
rect 460 -440 480 -380
rect 380 -460 480 -440
rect 520 -380 620 -360
rect 520 -440 540 -380
rect 600 -440 620 -380
rect 520 -460 620 -440
rect 660 -380 760 -360
rect 660 -440 680 -380
rect 740 -440 760 -380
rect 660 -460 760 -440
rect 800 -380 900 -360
rect 800 -440 820 -380
rect 880 -440 900 -380
rect 800 -460 900 -440
rect 940 -380 1040 -360
rect 940 -440 960 -380
rect 1020 -440 1040 -380
rect 940 -460 1040 -440
rect 1080 -380 1180 -360
rect 1080 -440 1100 -380
rect 1160 -440 1180 -380
rect 1080 -460 1180 -440
rect 1220 -380 1320 -360
rect 1220 -440 1240 -380
rect 1300 -440 1320 -380
rect 1220 -460 1320 -440
rect 4590 -510 5010 -490
rect 4590 -550 4950 -510
rect 4990 -550 5010 -510
rect 4590 -560 5010 -550
rect 4590 -620 4670 -560
rect 720 -720 820 -620
rect 4590 -660 4610 -620
rect 4650 -660 4670 -620
rect 4590 -790 4670 -660
rect 4710 -620 4770 -600
rect 4710 -660 4720 -620
rect 4760 -660 4770 -620
rect 4710 -690 4770 -660
rect 4900 -620 4960 -600
rect 4900 -660 4910 -620
rect 4950 -660 4960 -620
rect 4900 -690 4960 -660
rect 5090 -630 5150 -600
rect 5090 -670 5100 -630
rect 5140 -670 5150 -630
rect 5090 -690 5150 -670
rect 5190 -630 5270 -490
rect 5190 -670 5210 -630
rect 5250 -670 5270 -630
rect 5190 -730 5270 -670
rect 4850 -770 4870 -730
rect 4910 -770 5270 -730
rect 4850 -790 5270 -770
<< viali >>
rect 5590 -120 5630 -80
rect 5770 -120 5810 -80
rect 400 -280 460 -220
rect 203 -320 237 -286
rect 540 -280 600 -220
rect 680 -280 740 -220
rect 820 -280 880 -220
rect 960 -280 1020 -220
rect 1100 -280 1160 -220
rect 1240 -280 1300 -220
rect 60 -440 120 -380
rect 400 -440 460 -380
rect 540 -440 600 -380
rect 680 -440 740 -380
rect 820 -440 880 -380
rect 960 -440 1020 -380
rect 1100 -440 1160 -380
rect 1240 -440 1300 -380
rect 4610 -660 4650 -620
rect 4720 -660 4760 -620
rect 4910 -660 4950 -620
rect 5100 -670 5140 -630
rect 5210 -670 5250 -630
<< metal1 >>
rect 200 180 1800 220
rect 4420 160 4460 940
rect 4490 160 4520 940
rect 5310 210 5390 280
rect 5310 150 5320 210
rect 5380 150 5390 210
rect 5310 80 5390 150
rect 5570 -20 5690 10
rect 5580 -80 5640 -60
rect 5580 -120 5590 -80
rect 5630 -120 5640 -80
rect 5580 -140 5640 -120
rect 5760 -80 5820 -60
rect 5760 -120 5770 -80
rect 5810 -120 5820 -80
rect 5760 -140 5820 -120
rect 380 -220 480 -200
rect 380 -280 400 -220
rect 460 -280 480 -220
rect 191 -286 249 -280
rect 191 -320 203 -286
rect 237 -320 249 -286
rect 380 -300 480 -280
rect 520 -220 620 -140
rect 520 -280 540 -220
rect 600 -280 620 -220
rect 520 -300 620 -280
rect 660 -220 760 -200
rect 660 -280 680 -220
rect 740 -280 760 -220
rect 660 -300 760 -280
rect 800 -220 900 -200
rect 800 -280 820 -220
rect 880 -280 900 -220
rect 800 -300 900 -280
rect 940 -220 1040 -200
rect 940 -280 960 -220
rect 1020 -280 1040 -220
rect 940 -300 1040 -280
rect 1080 -220 1180 -200
rect 1080 -280 1100 -220
rect 1160 -280 1180 -220
rect 1080 -300 1180 -280
rect 1220 -220 1320 -200
rect 1220 -280 1240 -220
rect 1300 -280 1320 -220
rect 1220 -300 1320 -280
rect 191 -326 249 -320
rect 40 -380 140 -360
rect 40 -440 60 -380
rect 120 -440 140 -380
rect 40 -460 140 -440
rect 380 -380 480 -360
rect 380 -440 400 -380
rect 460 -440 480 -380
rect 380 -460 480 -440
rect 520 -380 620 -360
rect 520 -440 540 -380
rect 600 -440 620 -380
rect 520 -460 620 -440
rect 660 -380 760 -360
rect 660 -440 680 -380
rect 740 -440 760 -380
rect 660 -460 760 -440
rect 800 -380 900 -360
rect 800 -440 820 -380
rect 880 -440 900 -380
rect 800 -460 900 -440
rect 940 -380 1040 -360
rect 940 -440 960 -380
rect 1020 -440 1040 -380
rect 940 -460 1040 -440
rect 1080 -380 1180 -360
rect 1080 -440 1100 -380
rect 1160 -440 1180 -380
rect 1080 -460 1180 -440
rect 1220 -380 1320 -360
rect 1220 -440 1240 -380
rect 1300 -440 1320 -380
rect 1220 -460 1320 -440
rect 4590 -580 5310 -550
rect 4590 -620 4670 -610
rect 4720 -614 4760 -580
rect 900 -720 1000 -620
rect 4590 -660 4610 -620
rect 4650 -660 4670 -620
rect 4590 -670 4670 -660
rect 4708 -620 4772 -614
rect 4708 -660 4720 -620
rect 4760 -660 4772 -620
rect 4708 -666 4772 -660
rect 4890 -670 4900 -610
rect 4960 -670 4970 -610
rect 5088 -630 5152 -624
rect 5088 -670 5100 -630
rect 5140 -670 5152 -630
rect 5088 -676 5152 -670
rect 5190 -630 5270 -620
rect 5190 -670 5210 -630
rect 5250 -670 5270 -630
rect 5100 -710 5140 -676
rect 5190 -680 5270 -670
rect 4590 -740 5310 -710
<< via1 >>
rect 5320 150 5380 210
rect 540 -280 600 -220
rect 60 -440 120 -380
rect 4900 -620 4960 -610
rect 4900 -660 4910 -620
rect 4910 -660 4950 -620
rect 4950 -660 4960 -620
rect 4900 -670 4960 -660
<< metal2 >>
rect 5320 250 5430 280
rect 200 180 1800 220
rect 5320 210 5380 220
rect 5320 140 5380 150
rect 520 -220 620 -200
rect 520 -280 540 -220
rect 600 -280 620 -220
rect 520 -360 620 -280
rect 40 -380 140 -360
rect 40 -440 60 -380
rect 120 -440 140 -380
rect 40 -460 140 -440
rect 4900 -610 4960 -450
rect 1070 -720 1170 -620
rect 4900 -790 4960 -670
use dram3t_alpha  dram3t_alpha_0
timestamp 1719752019
transform -1 0 8112 0 -1 -1260
box 3920 -2120 4662 -1700
use dram3t_alpha  dram3t_alpha_1
timestamp 1719752019
transform -1 0 7652 0 -1 -1000
box 3920 -2120 4662 -1700
use dram3t_alpha  dram3t_alpha_2
timestamp 1719752019
transform -1 0 8112 0 -1 -1000
box 3920 -2120 4662 -1700
use dram3t_alpha  dram3t_alpha_3
timestamp 1719752019
transform -1 0 8112 0 -1 -1520
box 3920 -2120 4662 -1700
use dram3t_alpha  dram3t_alpha_4
timestamp 1719752019
transform -1 0 7652 0 -1 -1260
box 3920 -2120 4662 -1700
use dram3t_alpha  dram3t_alpha_5
timestamp 1719752019
transform -1 0 7652 0 -1 -1520
box 3920 -2120 4662 -1700
use dram3t_charlie  dram3t_charlie_0
array 0 2 720 0 5 340
timestamp 1719784265
transform 1 0 1030 0 1 1760
box -5270 -6820 -4550 -6460
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_0
timestamp 1719781273
transform 1 0 5738 0 1 -521
box -211 -252 211 252
<< labels >>
flabel locali 1760 -80 1800 -40 0 FreeSans 1600 0 0 0 C1N
flabel metal1 200 180 240 220 0 FreeSans 1600 0 0 0 C2M1
flabel metal2 1760 180 1800 220 0 FreeSans 1600 0 0 0 C2M2
flabel locali 258 -426 270 -386 0 FreeSans 800 90 32 0 TD
port 3 nsew
flabel locali 170 -412 182 -372 0 FreeSans 800 90 32 0 TS
port 5 nsew
flabel viali 203 -320 237 -286 0 FreeSans 800 0 0 0 TG
port 6 nsew
flabel locali 550 -300 580 -280 0 FreeSans 320 0 0 0 ARR_S
flabel locali 750 -690 820 -670 0 FreeSans 320 90 0 0 SINGLE_LI
flabel metal1 920 -680 960 -660 0 FreeSans 320 90 0 0 SINGLE_M1
flabel metal2 1100 -680 1140 -660 0 FreeSans 320 90 0 0 SINGLE_M2
flabel poly 550 -690 590 -650 0 FreeSans 320 0 0 0 SINGLE_P
flabel poly 200 -80 240 -40 0 FreeSans 1600 0 0 0 C1P
flabel poly 4890 300 4920 330 0 FreeSans 160 90 0 0 RD
flabel poly 4780 300 4810 330 0 FreeSans 160 90 0 0 WRB
flabel poly 5000 300 5030 330 0 FreeSans 160 90 0 0 SG
flabel ndiffc 4830 230 4870 270 0 FreeSans 320 90 0 0 BL
flabel ndiffc 4940 -60 4980 -20 0 FreeSans 320 90 0 0 BLB
flabel poly 5000 10 5030 40 0 FreeSans 160 90 0 0 WR
flabel poly 4780 10 4810 40 0 FreeSans 160 90 0 0 SGB
flabel poly 4890 10 4920 40 0 FreeSans 160 90 0 0 RDB
flabel ndiffc 4910 -660 4950 -620 0 FreeSans 160 90 0 0 VS
flabel ndiff 4730 -660 4770 -620 0 FreeSans 160 90 0 0 BL
flabel ndiff 5100 -660 5140 -620 0 FreeSans 160 90 0 0 BLB
flabel poly 5050 -500 5080 -470 0 FreeSans 160 90 0 0 RDB
flabel poly 4780 -770 4810 -740 0 FreeSans 160 90 0 0 RD
flabel poly 5160 -500 5190 -470 0 FreeSans 160 90 0 0 WR
flabel poly 4670 -770 4700 -740 0 FreeSans 160 90 0 0 WRB
flabel locali 4590 -530 4620 -500 0 FreeSans 160 90 0 0 VGB
flabel locali 5240 -770 5270 -740 0 FreeSans 160 90 0 0 VG
<< properties >>
string FIXED_BBOX -158 -199 158 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
