magic
tech sky130A
magscale 1 2
timestamp 1725372531
<< pwell >>
rect -1273 -567 1273 567
<< mvnmos >>
rect -1045 109 -845 309
rect -667 109 -467 309
rect -289 109 -89 309
rect 89 109 289 309
rect 467 109 667 309
rect 845 109 1045 309
rect -1045 -309 -845 -109
rect -667 -309 -467 -109
rect -289 -309 -89 -109
rect 89 -309 289 -109
rect 467 -309 667 -109
rect 845 -309 1045 -109
<< mvndiff >>
rect -1103 297 -1045 309
rect -1103 121 -1091 297
rect -1057 121 -1045 297
rect -1103 109 -1045 121
rect -845 297 -787 309
rect -845 121 -833 297
rect -799 121 -787 297
rect -845 109 -787 121
rect -725 297 -667 309
rect -725 121 -713 297
rect -679 121 -667 297
rect -725 109 -667 121
rect -467 297 -409 309
rect -467 121 -455 297
rect -421 121 -409 297
rect -467 109 -409 121
rect -347 297 -289 309
rect -347 121 -335 297
rect -301 121 -289 297
rect -347 109 -289 121
rect -89 297 -31 309
rect -89 121 -77 297
rect -43 121 -31 297
rect -89 109 -31 121
rect 31 297 89 309
rect 31 121 43 297
rect 77 121 89 297
rect 31 109 89 121
rect 289 297 347 309
rect 289 121 301 297
rect 335 121 347 297
rect 289 109 347 121
rect 409 297 467 309
rect 409 121 421 297
rect 455 121 467 297
rect 409 109 467 121
rect 667 297 725 309
rect 667 121 679 297
rect 713 121 725 297
rect 667 109 725 121
rect 787 297 845 309
rect 787 121 799 297
rect 833 121 845 297
rect 787 109 845 121
rect 1045 297 1103 309
rect 1045 121 1057 297
rect 1091 121 1103 297
rect 1045 109 1103 121
rect -1103 -121 -1045 -109
rect -1103 -297 -1091 -121
rect -1057 -297 -1045 -121
rect -1103 -309 -1045 -297
rect -845 -121 -787 -109
rect -845 -297 -833 -121
rect -799 -297 -787 -121
rect -845 -309 -787 -297
rect -725 -121 -667 -109
rect -725 -297 -713 -121
rect -679 -297 -667 -121
rect -725 -309 -667 -297
rect -467 -121 -409 -109
rect -467 -297 -455 -121
rect -421 -297 -409 -121
rect -467 -309 -409 -297
rect -347 -121 -289 -109
rect -347 -297 -335 -121
rect -301 -297 -289 -121
rect -347 -309 -289 -297
rect -89 -121 -31 -109
rect -89 -297 -77 -121
rect -43 -297 -31 -121
rect -89 -309 -31 -297
rect 31 -121 89 -109
rect 31 -297 43 -121
rect 77 -297 89 -121
rect 31 -309 89 -297
rect 289 -121 347 -109
rect 289 -297 301 -121
rect 335 -297 347 -121
rect 289 -309 347 -297
rect 409 -121 467 -109
rect 409 -297 421 -121
rect 455 -297 467 -121
rect 409 -309 467 -297
rect 667 -121 725 -109
rect 667 -297 679 -121
rect 713 -297 725 -121
rect 667 -309 725 -297
rect 787 -121 845 -109
rect 787 -297 799 -121
rect 833 -297 845 -121
rect 787 -309 845 -297
rect 1045 -121 1103 -109
rect 1045 -297 1057 -121
rect 1091 -297 1103 -121
rect 1045 -309 1103 -297
<< mvndiffc >>
rect -1091 121 -1057 297
rect -833 121 -799 297
rect -713 121 -679 297
rect -455 121 -421 297
rect -335 121 -301 297
rect -77 121 -43 297
rect 43 121 77 297
rect 301 121 335 297
rect 421 121 455 297
rect 679 121 713 297
rect 799 121 833 297
rect 1057 121 1091 297
rect -1091 -297 -1057 -121
rect -833 -297 -799 -121
rect -713 -297 -679 -121
rect -455 -297 -421 -121
rect -335 -297 -301 -121
rect -77 -297 -43 -121
rect 43 -297 77 -121
rect 301 -297 335 -121
rect 421 -297 455 -121
rect 679 -297 713 -121
rect 799 -297 833 -121
rect 1057 -297 1091 -121
<< mvpsubdiff >>
rect -1237 519 1237 531
rect -1237 485 -1129 519
rect 1129 485 1237 519
rect -1237 473 1237 485
rect -1237 423 -1179 473
rect -1237 -423 -1225 423
rect -1191 -423 -1179 423
rect 1179 423 1237 473
rect -1237 -473 -1179 -423
rect 1179 -423 1191 423
rect 1225 -423 1237 423
rect 1179 -473 1237 -423
rect -1237 -485 1237 -473
rect -1237 -519 -1129 -485
rect 1129 -519 1237 -485
rect -1237 -531 1237 -519
<< mvpsubdiffcont >>
rect -1129 485 1129 519
rect -1225 -423 -1191 423
rect 1191 -423 1225 423
rect -1129 -519 1129 -485
<< poly >>
rect -1045 381 -845 397
rect -1045 347 -1029 381
rect -861 347 -845 381
rect -1045 309 -845 347
rect -667 381 -467 397
rect -667 347 -651 381
rect -483 347 -467 381
rect -667 309 -467 347
rect -289 381 -89 397
rect -289 347 -273 381
rect -105 347 -89 381
rect -289 309 -89 347
rect 89 381 289 397
rect 89 347 105 381
rect 273 347 289 381
rect 89 309 289 347
rect 467 381 667 397
rect 467 347 483 381
rect 651 347 667 381
rect 467 309 667 347
rect 845 381 1045 397
rect 845 347 861 381
rect 1029 347 1045 381
rect 845 309 1045 347
rect -1045 71 -845 109
rect -1045 37 -1029 71
rect -861 37 -845 71
rect -1045 21 -845 37
rect -667 71 -467 109
rect -667 37 -651 71
rect -483 37 -467 71
rect -667 21 -467 37
rect -289 71 -89 109
rect -289 37 -273 71
rect -105 37 -89 71
rect -289 21 -89 37
rect 89 71 289 109
rect 89 37 105 71
rect 273 37 289 71
rect 89 21 289 37
rect 467 71 667 109
rect 467 37 483 71
rect 651 37 667 71
rect 467 21 667 37
rect 845 71 1045 109
rect 845 37 861 71
rect 1029 37 1045 71
rect 845 21 1045 37
rect -1045 -37 -845 -21
rect -1045 -71 -1029 -37
rect -861 -71 -845 -37
rect -1045 -109 -845 -71
rect -667 -37 -467 -21
rect -667 -71 -651 -37
rect -483 -71 -467 -37
rect -667 -109 -467 -71
rect -289 -37 -89 -21
rect -289 -71 -273 -37
rect -105 -71 -89 -37
rect -289 -109 -89 -71
rect 89 -37 289 -21
rect 89 -71 105 -37
rect 273 -71 289 -37
rect 89 -109 289 -71
rect 467 -37 667 -21
rect 467 -71 483 -37
rect 651 -71 667 -37
rect 467 -109 667 -71
rect 845 -37 1045 -21
rect 845 -71 861 -37
rect 1029 -71 1045 -37
rect 845 -109 1045 -71
rect -1045 -347 -845 -309
rect -1045 -381 -1029 -347
rect -861 -381 -845 -347
rect -1045 -397 -845 -381
rect -667 -347 -467 -309
rect -667 -381 -651 -347
rect -483 -381 -467 -347
rect -667 -397 -467 -381
rect -289 -347 -89 -309
rect -289 -381 -273 -347
rect -105 -381 -89 -347
rect -289 -397 -89 -381
rect 89 -347 289 -309
rect 89 -381 105 -347
rect 273 -381 289 -347
rect 89 -397 289 -381
rect 467 -347 667 -309
rect 467 -381 483 -347
rect 651 -381 667 -347
rect 467 -397 667 -381
rect 845 -347 1045 -309
rect 845 -381 861 -347
rect 1029 -381 1045 -347
rect 845 -397 1045 -381
<< polycont >>
rect -1029 347 -861 381
rect -651 347 -483 381
rect -273 347 -105 381
rect 105 347 273 381
rect 483 347 651 381
rect 861 347 1029 381
rect -1029 37 -861 71
rect -651 37 -483 71
rect -273 37 -105 71
rect 105 37 273 71
rect 483 37 651 71
rect 861 37 1029 71
rect -1029 -71 -861 -37
rect -651 -71 -483 -37
rect -273 -71 -105 -37
rect 105 -71 273 -37
rect 483 -71 651 -37
rect 861 -71 1029 -37
rect -1029 -381 -861 -347
rect -651 -381 -483 -347
rect -273 -381 -105 -347
rect 105 -381 273 -347
rect 483 -381 651 -347
rect 861 -381 1029 -347
<< locali >>
rect -1225 485 -1129 519
rect 1129 485 1225 519
rect -1225 423 -1191 485
rect 1191 423 1225 485
rect -1045 347 -1029 381
rect -861 347 -845 381
rect -667 347 -651 381
rect -483 347 -467 381
rect -289 347 -273 381
rect -105 347 -89 381
rect 89 347 105 381
rect 273 347 289 381
rect 467 347 483 381
rect 651 347 667 381
rect 845 347 861 381
rect 1029 347 1045 381
rect -1091 297 -1057 313
rect -1091 105 -1057 121
rect -833 297 -799 313
rect -833 105 -799 121
rect -713 297 -679 313
rect -713 105 -679 121
rect -455 297 -421 313
rect -455 105 -421 121
rect -335 297 -301 313
rect -335 105 -301 121
rect -77 297 -43 313
rect -77 105 -43 121
rect 43 297 77 313
rect 43 105 77 121
rect 301 297 335 313
rect 301 105 335 121
rect 421 297 455 313
rect 421 105 455 121
rect 679 297 713 313
rect 679 105 713 121
rect 799 297 833 313
rect 799 105 833 121
rect 1057 297 1091 313
rect 1057 105 1091 121
rect -1045 37 -1029 71
rect -861 37 -845 71
rect -667 37 -651 71
rect -483 37 -467 71
rect -289 37 -273 71
rect -105 37 -89 71
rect 89 37 105 71
rect 273 37 289 71
rect 467 37 483 71
rect 651 37 667 71
rect 845 37 861 71
rect 1029 37 1045 71
rect -1045 -71 -1029 -37
rect -861 -71 -845 -37
rect -667 -71 -651 -37
rect -483 -71 -467 -37
rect -289 -71 -273 -37
rect -105 -71 -89 -37
rect 89 -71 105 -37
rect 273 -71 289 -37
rect 467 -71 483 -37
rect 651 -71 667 -37
rect 845 -71 861 -37
rect 1029 -71 1045 -37
rect -1091 -121 -1057 -105
rect -1091 -313 -1057 -297
rect -833 -121 -799 -105
rect -833 -313 -799 -297
rect -713 -121 -679 -105
rect -713 -313 -679 -297
rect -455 -121 -421 -105
rect -455 -313 -421 -297
rect -335 -121 -301 -105
rect -335 -313 -301 -297
rect -77 -121 -43 -105
rect -77 -313 -43 -297
rect 43 -121 77 -105
rect 43 -313 77 -297
rect 301 -121 335 -105
rect 301 -313 335 -297
rect 421 -121 455 -105
rect 421 -313 455 -297
rect 679 -121 713 -105
rect 679 -313 713 -297
rect 799 -121 833 -105
rect 799 -313 833 -297
rect 1057 -121 1091 -105
rect 1057 -313 1091 -297
rect -1045 -381 -1029 -347
rect -861 -381 -845 -347
rect -667 -381 -651 -347
rect -483 -381 -467 -347
rect -289 -381 -273 -347
rect -105 -381 -89 -347
rect 89 -381 105 -347
rect 273 -381 289 -347
rect 467 -381 483 -347
rect 651 -381 667 -347
rect 845 -381 861 -347
rect 1029 -381 1045 -347
rect -1225 -485 -1191 -423
rect 1191 -485 1225 -423
rect -1225 -519 -1129 -485
rect 1129 -519 1225 -485
<< viali >>
rect -1225 -388 -1191 388
rect -1029 347 -861 381
rect -651 347 -483 381
rect -273 347 -105 381
rect 105 347 273 381
rect 483 347 651 381
rect 861 347 1029 381
rect -1091 138 -1057 208
rect -833 210 -799 280
rect -713 210 -679 280
rect -455 138 -421 208
rect -335 138 -301 208
rect -77 210 -43 280
rect 43 210 77 280
rect 301 138 335 208
rect 421 138 455 208
rect 679 210 713 280
rect 799 210 833 280
rect 1057 138 1091 208
rect -1029 37 -861 71
rect -651 37 -483 71
rect -273 37 -105 71
rect 105 37 273 71
rect 483 37 651 71
rect 861 37 1029 71
rect -1029 -71 -861 -37
rect -651 -71 -483 -37
rect -273 -71 -105 -37
rect 105 -71 273 -37
rect 483 -71 651 -37
rect 861 -71 1029 -37
rect -1091 -280 -1057 -210
rect -833 -208 -799 -138
rect -713 -208 -679 -138
rect -455 -280 -421 -210
rect -335 -280 -301 -210
rect -77 -208 -43 -138
rect 43 -208 77 -138
rect 301 -280 335 -210
rect 421 -280 455 -210
rect 679 -208 713 -138
rect 799 -208 833 -138
rect 1057 -280 1091 -210
rect -1029 -381 -861 -347
rect -651 -381 -483 -347
rect -273 -381 -105 -347
rect 105 -381 273 -347
rect 483 -381 651 -347
rect 861 -381 1029 -347
rect 1191 -388 1225 388
rect -953 -519 953 -485
<< metal1 >>
rect -1231 388 -1185 400
rect -1231 -388 -1225 388
rect -1191 -388 -1185 388
rect 1185 388 1231 400
rect -1041 381 -849 387
rect -1041 347 -1029 381
rect -861 347 -849 381
rect -1041 341 -849 347
rect -663 381 -471 387
rect -663 347 -651 381
rect -483 347 -471 381
rect -663 341 -471 347
rect -285 381 -93 387
rect -285 347 -273 381
rect -105 347 -93 381
rect -285 341 -93 347
rect 93 381 285 387
rect 93 347 105 381
rect 273 347 285 381
rect 93 341 285 347
rect 471 381 663 387
rect 471 347 483 381
rect 651 347 663 381
rect 471 341 663 347
rect 849 381 1041 387
rect 849 347 861 381
rect 1029 347 1041 381
rect 849 341 1041 347
rect -839 280 -793 292
rect -1097 208 -1051 220
rect -1097 138 -1091 208
rect -1057 138 -1051 208
rect -839 210 -833 280
rect -799 210 -793 280
rect -839 198 -793 210
rect -719 280 -673 292
rect -719 210 -713 280
rect -679 210 -673 280
rect -83 280 -37 292
rect -719 198 -673 210
rect -461 208 -415 220
rect -1097 126 -1051 138
rect -461 138 -455 208
rect -421 138 -415 208
rect -461 126 -415 138
rect -341 208 -295 220
rect -341 138 -335 208
rect -301 138 -295 208
rect -83 210 -77 280
rect -43 210 -37 280
rect -83 198 -37 210
rect 37 280 83 292
rect 37 210 43 280
rect 77 210 83 280
rect 673 280 719 292
rect 37 198 83 210
rect 295 208 341 220
rect -341 126 -295 138
rect 295 138 301 208
rect 335 138 341 208
rect 295 126 341 138
rect 415 208 461 220
rect 415 138 421 208
rect 455 138 461 208
rect 673 210 679 280
rect 713 210 719 280
rect 673 198 719 210
rect 793 280 839 292
rect 793 210 799 280
rect 833 210 839 280
rect 793 198 839 210
rect 1051 208 1097 220
rect 415 126 461 138
rect 1051 138 1057 208
rect 1091 138 1097 208
rect 1051 126 1097 138
rect -1041 71 -849 77
rect -1041 37 -1029 71
rect -861 37 -849 71
rect -1041 31 -849 37
rect -663 71 -471 77
rect -663 37 -651 71
rect -483 37 -471 71
rect -663 31 -471 37
rect -285 71 -93 77
rect -285 37 -273 71
rect -105 37 -93 71
rect -285 31 -93 37
rect 93 71 285 77
rect 93 37 105 71
rect 273 37 285 71
rect 93 31 285 37
rect 471 71 663 77
rect 471 37 483 71
rect 651 37 663 71
rect 471 31 663 37
rect 849 71 1041 77
rect 849 37 861 71
rect 1029 37 1041 71
rect 849 31 1041 37
rect -1041 -37 -849 -31
rect -1041 -71 -1029 -37
rect -861 -71 -849 -37
rect -1041 -77 -849 -71
rect -663 -37 -471 -31
rect -663 -71 -651 -37
rect -483 -71 -471 -37
rect -663 -77 -471 -71
rect -285 -37 -93 -31
rect -285 -71 -273 -37
rect -105 -71 -93 -37
rect -285 -77 -93 -71
rect 93 -37 285 -31
rect 93 -71 105 -37
rect 273 -71 285 -37
rect 93 -77 285 -71
rect 471 -37 663 -31
rect 471 -71 483 -37
rect 651 -71 663 -37
rect 471 -77 663 -71
rect 849 -37 1041 -31
rect 849 -71 861 -37
rect 1029 -71 1041 -37
rect 849 -77 1041 -71
rect -839 -138 -793 -126
rect -1097 -210 -1051 -198
rect -1097 -280 -1091 -210
rect -1057 -280 -1051 -210
rect -839 -208 -833 -138
rect -799 -208 -793 -138
rect -839 -220 -793 -208
rect -719 -138 -673 -126
rect -719 -208 -713 -138
rect -679 -208 -673 -138
rect -83 -138 -37 -126
rect -719 -220 -673 -208
rect -461 -210 -415 -198
rect -1097 -292 -1051 -280
rect -461 -280 -455 -210
rect -421 -280 -415 -210
rect -461 -292 -415 -280
rect -341 -210 -295 -198
rect -341 -280 -335 -210
rect -301 -280 -295 -210
rect -83 -208 -77 -138
rect -43 -208 -37 -138
rect -83 -220 -37 -208
rect 37 -138 83 -126
rect 37 -208 43 -138
rect 77 -208 83 -138
rect 673 -138 719 -126
rect 37 -220 83 -208
rect 295 -210 341 -198
rect -341 -292 -295 -280
rect 295 -280 301 -210
rect 335 -280 341 -210
rect 295 -292 341 -280
rect 415 -210 461 -198
rect 415 -280 421 -210
rect 455 -280 461 -210
rect 673 -208 679 -138
rect 713 -208 719 -138
rect 673 -220 719 -208
rect 793 -138 839 -126
rect 793 -208 799 -138
rect 833 -208 839 -138
rect 793 -220 839 -208
rect 1051 -210 1097 -198
rect 415 -292 461 -280
rect 1051 -280 1057 -210
rect 1091 -280 1097 -210
rect 1051 -292 1097 -280
rect -1041 -347 -849 -341
rect -1041 -381 -1029 -347
rect -861 -381 -849 -347
rect -1041 -387 -849 -381
rect -663 -347 -471 -341
rect -663 -381 -651 -347
rect -483 -381 -471 -347
rect -663 -387 -471 -381
rect -285 -347 -93 -341
rect -285 -381 -273 -347
rect -105 -381 -93 -347
rect -285 -387 -93 -381
rect 93 -347 285 -341
rect 93 -381 105 -347
rect 273 -381 285 -347
rect 93 -387 285 -381
rect 471 -347 663 -341
rect 471 -381 483 -347
rect 651 -381 663 -347
rect 471 -387 663 -381
rect 849 -347 1041 -341
rect 849 -381 861 -347
rect 1029 -381 1041 -347
rect 849 -387 1041 -381
rect -1231 -400 -1185 -388
rect 1185 -388 1191 388
rect 1225 -388 1231 388
rect 1185 -400 1231 -388
rect -965 -485 965 -479
rect -965 -519 -953 -485
rect 953 -519 965 -485
rect -965 -525 965 -519
<< properties >>
string FIXED_BBOX -1208 -502 1208 502
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 2 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 80 viagr 80 viagl 80 viagt 0
string sky130_fd_pr__nfet_g5v0d10v5_HF5BS6 parameters
<< end >>
