magic
tech sky130A
magscale 1 2
timestamp 1725372531
<< pwell >>
rect -2120 -200 -1980 -100
<< locali >>
rect -3040 1660 320 1720
rect -3040 1560 -2700 1660
rect 120 1560 320 1660
rect -3040 1440 320 1560
rect -3040 440 -2920 1440
rect -3040 360 -3020 440
rect -2940 420 -2920 440
rect -2940 360 -2340 420
rect -2260 360 -1780 420
rect 200 420 320 1440
rect -1700 360 -280 420
rect -3040 340 -280 360
rect -200 340 220 420
rect 300 340 320 420
rect -3040 320 320 340
rect -3040 60 320 100
rect -3040 -20 -2660 60
rect -3040 -1040 -2940 -20
rect -2780 -1040 -2660 -20
rect -2460 40 320 60
rect -100 -20 320 40
rect -100 -940 60 -20
rect -2460 -1020 -2420 -940
rect -140 -1020 60 -940
rect -2460 -1040 60 -1020
rect 220 -1040 320 -20
rect -3040 -1080 320 -1040
<< viali >>
rect -2700 1560 120 1660
rect -3020 360 -2940 440
rect -2340 360 -2260 440
rect -1780 360 -1700 440
rect -280 340 -200 420
rect 220 340 300 420
rect -2940 -1040 -2780 -20
rect -2660 -1040 -2460 60
rect -2420 -1020 -140 -940
rect 60 -1040 220 -20
<< metal1 >>
rect -3040 1660 320 1720
rect -3040 1560 -2700 1660
rect 120 1560 320 1660
rect -3040 1510 320 1560
rect -3040 1430 -2920 1510
rect -2840 1430 320 1510
rect -3040 1400 320 1430
rect -3040 1060 -2830 1400
rect -2720 1070 -2660 1340
rect -2570 1210 -2420 1260
rect -2570 1090 -2550 1210
rect -2430 1090 -2420 1210
rect -3040 440 -2920 1060
rect -2750 1010 -2740 1070
rect -2780 970 -2740 1010
rect -2640 1010 -2630 1070
rect -2570 1050 -2420 1090
rect -2330 1010 -2270 1340
rect -2180 1060 -2060 1400
rect -1950 1010 -1890 1340
rect -1810 1210 -1660 1260
rect -1810 1090 -1800 1210
rect -1680 1090 -1660 1210
rect -1810 1050 -1660 1090
rect -1580 1010 -1520 1340
rect -1420 1050 -1300 1400
rect -1200 1010 -1140 1340
rect -1060 1210 -900 1260
rect -1060 1090 -1050 1210
rect -930 1090 -900 1210
rect -1060 1070 -900 1090
rect -820 1010 -760 1340
rect -660 1050 -540 1400
rect -460 1010 -400 1340
rect -310 1210 -150 1250
rect -310 1090 -290 1210
rect -170 1090 -150 1210
rect -310 1060 -150 1090
rect -60 1040 0 1340
rect 90 1060 320 1400
rect -90 1010 -80 1040
rect -2640 970 -1450 1010
rect -2780 960 -1450 970
rect -1260 960 -80 1010
rect 0 1010 10 1040
rect 0 960 70 1010
rect -2840 860 90 920
rect -2840 610 -2690 860
rect -2570 770 -2420 820
rect -2570 650 -2550 770
rect -2430 650 -2420 770
rect -2570 610 -2420 650
rect -2300 610 -2150 860
rect -2110 610 -1960 860
rect -1810 770 -1660 820
rect -1810 650 -1800 770
rect -1680 650 -1660 770
rect -1810 610 -1660 650
rect -1510 610 -1390 860
rect -1350 650 -1340 770
rect -1260 650 -1250 770
rect -2750 530 -2690 610
rect -2300 540 -2240 610
rect -2020 540 -1960 610
rect -1510 540 -1400 610
rect -1200 540 -1140 860
rect -1060 780 -900 820
rect -1060 660 -1050 780
rect -930 660 -900 780
rect -1060 640 -900 660
rect -2352 440 -2248 446
rect -1792 440 -1688 446
rect -3040 360 -3020 440
rect -2940 360 -2340 440
rect -2260 360 -1780 440
rect -1700 360 -1600 440
rect -3040 340 -1600 360
rect -3040 250 -2960 260
rect -3040 170 -2010 250
rect -3040 160 -2960 170
rect -2666 60 -2454 72
rect -3040 -20 -2660 60
rect -3040 -1040 -2940 -20
rect -2780 -80 -2660 -20
rect -2780 -180 -2740 -80
rect -2780 -1040 -2660 -180
rect -2460 -920 -2454 60
rect -2090 -80 -2010 170
rect -1480 190 -1400 540
rect -820 530 -760 860
rect -680 620 -520 820
rect -660 600 -530 620
rect -630 360 -550 600
rect -460 530 -400 860
rect -310 780 -150 820
rect -310 660 -290 780
rect -170 660 -150 780
rect -310 640 -150 660
rect -60 540 0 860
rect 40 640 50 760
rect 130 640 140 760
rect -292 420 -188 426
rect 180 420 320 1060
rect -690 340 -490 360
rect -690 190 -670 340
rect -510 190 -490 340
rect -380 340 -280 420
rect -200 340 220 420
rect 300 340 320 420
rect -380 320 320 340
rect -1480 110 -1250 190
rect -690 160 -490 190
rect -2320 -140 -1780 -80
rect -2410 -340 -2400 -240
rect -2320 -340 -2310 -240
rect -2120 -380 -1980 -140
rect -1790 -340 -1780 -240
rect -1700 -340 -1690 -240
rect -1640 -340 -1630 -240
rect -1550 -340 -1540 -240
rect -2300 -400 -1780 -380
rect -1480 -400 -1420 -90
rect -1330 -160 -1250 110
rect -1350 -370 -1230 -160
rect -1150 -400 -1090 -90
rect -1040 -340 -1030 -240
rect -950 -340 -940 -240
rect -880 -340 -870 -240
rect -790 -340 -780 -240
rect -720 -400 -660 -90
rect -570 -160 -490 160
rect -100 -20 320 100
rect -590 -370 -470 -160
rect -390 -400 -330 -90
rect -280 -340 -270 -240
rect -190 -340 -180 -240
rect -2300 -440 -240 -400
rect -2320 -510 -1780 -500
rect -2320 -560 -2280 -510
rect -2290 -590 -2280 -560
rect -2200 -560 -1000 -510
rect -820 -520 -240 -510
rect -820 -560 -380 -520
rect -2200 -590 -2180 -560
rect -2290 -600 -2180 -590
rect -2410 -780 -2400 -680
rect -2320 -780 -2310 -680
rect -2240 -820 -2180 -600
rect -2320 -880 -2140 -820
rect -2100 -920 -1990 -600
rect -1900 -820 -1840 -560
rect -1790 -780 -1780 -680
rect -1700 -780 -1690 -680
rect -1640 -780 -1630 -680
rect -1550 -780 -1540 -680
rect -1960 -880 -1780 -820
rect -1480 -860 -1420 -560
rect -1340 -920 -1230 -600
rect -1150 -850 -1090 -560
rect -1040 -780 -1030 -680
rect -950 -780 -940 -680
rect -880 -780 -870 -680
rect -790 -780 -780 -680
rect -710 -850 -650 -560
rect -400 -600 -380 -560
rect -300 -560 -240 -520
rect -300 -600 -290 -560
rect -590 -920 -480 -600
rect -400 -850 -340 -600
rect -280 -780 -270 -680
rect -190 -780 -180 -680
rect -100 -920 60 -20
rect -2460 -940 60 -920
rect -2460 -1020 -2420 -940
rect -140 -1020 60 -940
rect -2460 -1040 60 -1020
rect 220 -1040 320 -20
rect -3040 -1080 320 -1040
<< via1 >>
rect -2920 1430 -2840 1510
rect -2550 1090 -2430 1210
rect -2740 970 -2640 1070
rect -1800 1090 -1680 1210
rect -1050 1090 -930 1210
rect -290 1090 -170 1210
rect -80 960 0 1040
rect -2550 650 -2430 770
rect -1800 650 -1680 770
rect -1340 650 -1260 770
rect -1050 660 -930 780
rect -2740 -180 -2660 -80
rect -2660 -180 -2640 -80
rect -290 660 -170 780
rect 50 640 130 760
rect -670 190 -510 340
rect -2400 -340 -2320 -240
rect -1780 -340 -1700 -240
rect -1630 -340 -1550 -240
rect -1030 -340 -950 -240
rect -870 -340 -790 -240
rect -270 -340 -190 -240
rect -2280 -590 -2200 -510
rect -2400 -780 -2320 -680
rect -1780 -780 -1700 -680
rect -1630 -780 -1550 -680
rect -1030 -780 -950 -680
rect -870 -780 -790 -680
rect -380 -600 -300 -520
rect -270 -780 -190 -680
<< metal2 >>
rect -2920 1510 -2840 1560
rect -2920 -510 -2840 1430
rect -2550 1210 -2430 1220
rect -1800 1210 -1680 1220
rect -2430 1090 -1800 1210
rect -2740 1070 -2640 1080
rect -2740 -80 -2640 970
rect -2550 770 -2430 1090
rect -1800 1080 -1680 1090
rect -1050 1210 -930 1220
rect -290 1210 -170 1220
rect -930 1090 -290 1210
rect -1050 780 -930 1090
rect -290 1080 -170 1090
rect -80 1040 0 1050
rect 0 960 320 1040
rect -80 950 0 960
rect -290 780 -170 790
rect -1800 770 -1680 780
rect -2430 650 -1800 770
rect -2550 640 -2430 650
rect -1800 640 -1680 650
rect -1340 770 -1260 780
rect -930 660 -290 780
rect -1050 650 -930 660
rect -290 650 -170 660
rect 50 760 130 770
rect -1340 300 -1260 650
rect -690 340 -490 360
rect -690 300 -670 340
rect -1340 220 -670 300
rect -690 190 -670 220
rect -510 300 -490 340
rect 50 320 130 640
rect 30 300 130 320
rect -510 220 130 300
rect -510 190 -490 220
rect -690 160 -490 190
rect -2740 -186 -2640 -180
rect -2400 -240 -2320 -230
rect -1780 -240 -1700 -230
rect -2410 -340 -2400 -240
rect -2320 -340 -1780 -240
rect -2400 -350 -2320 -340
rect -2280 -510 -2200 -500
rect -2920 -590 -2280 -510
rect -2280 -600 -2200 -590
rect -2400 -680 -2320 -670
rect -1780 -680 -1700 -340
rect -1630 -240 -1550 -230
rect -1030 -240 -950 -230
rect -1550 -340 -1030 -240
rect -1630 -350 -1550 -340
rect -2320 -780 -1780 -680
rect -2400 -790 -2320 -780
rect -1780 -790 -1700 -780
rect -1630 -680 -1550 -670
rect -1030 -680 -950 -340
rect -1550 -780 -1030 -680
rect -1630 -790 -1550 -780
rect -1030 -790 -950 -780
rect -870 -240 -790 -230
rect -270 -240 -190 -230
rect -790 -340 -270 -240
rect -870 -680 -790 -340
rect -270 -350 -190 -340
rect -380 -520 -300 -510
rect -300 -600 320 -520
rect -380 -610 -300 -600
rect -270 -680 -190 -670
rect -790 -780 -270 -680
rect -870 -790 -790 -780
rect -270 -790 -190 -780
use sky130_fd_pr__nfet_g5v0d10v5_HF5BS6  sky130_fd_pr__nfet_g5v0d10v5_HF5BS6_0
timestamp 1725372531
transform 1 0 -1287 0 1 -473
box -1273 -567 1273 567
use sky130_fd_pr__pfet_g5v0d10v5_U7XX7W  sky130_fd_pr__pfet_g5v0d10v5_U7XX7W_0
timestamp 1725372531
transform 1 0 -1359 0 1 935
box -1681 -615 1681 615
<< labels >>
flabel metal2 30 220 130 320 0 FreeSans 1280 0 0 0 VOUT
port 1 nsew
flabel metal1 -2980 -1000 -2780 -800 0 FreeSans 1280 0 0 0 VSS
port 2 nsew
flabel metal1 -3000 1500 -2800 1700 0 FreeSans 1280 0 0 0 VDD
port 3 nsew
flabel metal1 -3040 160 -2960 260 0 FreeSans 1280 0 0 0 IREF
port 4 nsew
flabel metal2 240 -600 320 -520 0 FreeSans 1280 0 0 0 DN
port 5 nsew
flabel metal2 240 960 320 1040 0 FreeSans 1280 0 0 0 UPB
port 6 nsew
<< end >>
