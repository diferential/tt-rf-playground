magic
tech sky130A
magscale 1 2
timestamp 1723344990
<< metal1 >>
rect -100 1020 500 1120
rect 160 900 240 1020
rect 30 780 40 840
rect 100 820 110 840
rect 100 780 340 820
rect 0 680 140 720
rect -100 540 -40 560
rect 0 540 40 680
rect -100 500 40 540
rect 0 120 40 500
rect 80 500 100 560
rect 160 500 170 560
rect 80 160 120 500
rect 260 460 300 720
rect 250 400 260 460
rect 320 400 330 460
rect 260 300 300 400
rect 200 160 240 260
rect 0 80 200 120
rect 320 40 440 260
rect -100 -60 500 40
<< via1 >>
rect 40 780 100 840
rect 100 500 160 560
rect 260 400 320 460
<< metal2 >>
rect 40 840 100 850
rect 100 780 140 840
rect 40 770 140 780
rect 100 570 140 770
rect 100 560 160 570
rect 160 500 480 540
rect 100 490 160 500
rect 420 480 480 500
rect 260 460 320 470
rect -100 400 260 440
rect -100 380 -40 400
rect 260 390 320 400
use sky130_fd_pr__nfet_01v8_lvt_ZDUAWA  sky130_fd_pr__nfet_01v8_lvt_ZDUAWA_0
timestamp 1723344990
transform 1 0 222 0 1 207
box -275 -260 275 260
use sky130_fd_pr__pfet_01v8_lvt_UT4KY6  sky130_fd_pr__pfet_01v8_lvt_UT4KY6_0
timestamp 1723344990
transform 1 0 192 0 1 831
box -295 -284 295 284
<< labels >>
flabel metal1 -100 500 -40 560 0 FreeSans 800 0 0 0 A
port 0 nsew
flabel metal2 -100 380 -40 440 0 FreeSans 800 0 0 0 B
port 1 nsew
flabel metal2 420 480 480 540 0 FreeSans 800 0 0 0 Q
port 2 nsew
flabel metal1 -100 1020 0 1120 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal1 -60 -60 40 40 0 FreeSans 800 0 0 0 VSS
port 4 nsew
<< end >>
