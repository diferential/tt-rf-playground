magic
tech sky130A
magscale 1 2
timestamp 1717260631
<< metal1 >>
rect 19720 41630 19900 41660
rect 19720 41550 19771 41630
rect 19851 41550 19900 41630
rect 19720 41530 19900 41550
rect 19611 41380 19691 41386
rect 16600 41110 16740 41116
rect 16740 40970 18171 41110
rect 19611 41000 19691 41300
rect 19771 41000 19851 41530
rect 16600 40964 16740 40970
<< via1 >>
rect 19771 41550 19851 41630
rect 19611 41300 19691 41380
rect 16600 40970 16740 41110
<< metal2 >>
rect 25530 43608 25630 43630
rect 25530 43552 25562 43608
rect 25618 43552 25630 43608
rect 25330 42018 25430 43170
rect 25330 41962 25342 42018
rect 25398 41962 25430 42018
rect 19720 41630 19900 41660
rect 19720 41550 19771 41630
rect 19851 41550 19900 41630
rect 19720 41530 19900 41550
rect 19590 41380 19710 41420
rect 19590 41300 19611 41380
rect 19691 41300 19710 41380
rect 24390 41368 24450 41640
rect 24700 41498 24760 41690
rect 24900 41658 24960 41840
rect 25100 41838 25160 41950
rect 25330 41890 25430 41962
rect 25100 41782 25102 41838
rect 25158 41782 25160 41838
rect 25530 41830 25630 43552
rect 25730 42298 25830 43160
rect 25730 42242 25762 42298
rect 25818 42242 25830 42298
rect 25730 41900 25830 42242
rect 25950 42638 26050 43150
rect 25950 42582 25982 42638
rect 26038 42582 26050 42638
rect 25950 41914 26050 42582
rect 25100 41780 25160 41782
rect 25102 41773 25158 41780
rect 24900 41602 24902 41658
rect 24958 41602 24960 41658
rect 24900 41600 24960 41602
rect 24902 41593 24958 41600
rect 24693 41442 24702 41498
rect 24758 41442 24767 41498
rect 24700 41440 24760 41442
rect 24390 41312 24392 41368
rect 24448 41312 24450 41368
rect 24390 41310 24450 41312
rect 24392 41303 24448 41310
rect 19590 41290 19710 41300
rect 16594 40970 16600 41110
rect 16740 40970 16746 41110
rect 16600 28215 17200 40970
rect 25380 28220 25980 29838
rect 16596 27625 16605 28215
rect 17195 27625 17204 28215
rect 16600 27620 17200 27625
rect 25380 27611 25980 27620
rect 28275 8895 28385 8904
rect 28275 8776 28385 8785
rect 20431 7600 20440 7800
rect 20640 7600 21230 7800
rect 19990 7300 20130 7500
rect 20330 7300 21220 7500
rect 19650 4300 21320 4600
rect 19650 1000 19950 4300
rect 20240 3700 21310 4000
rect 20240 1530 20540 3700
rect 20240 1221 20540 1230
rect 19530 970 20000 1000
rect 19530 670 19650 970
rect 19950 670 20000 970
rect 19530 620 20000 670
<< via2 >>
rect 25562 43552 25618 43608
rect 25342 41962 25398 42018
rect 19771 41550 19851 41630
rect 19611 41300 19691 41380
rect 25102 41782 25158 41838
rect 25762 42242 25818 42298
rect 25982 42582 26038 42638
rect 24902 41602 24958 41658
rect 24702 41442 24758 41498
rect 24392 41312 24448 41368
rect 16605 27625 17195 28215
rect 25380 27620 25980 28220
rect 28275 8785 28385 8895
rect 20440 7600 20640 7800
rect 20130 7300 20330 7500
rect 20240 1230 20540 1530
rect 19650 670 19950 970
<< metal3 >>
rect 20130 43899 23210 43900
rect 20125 43701 20131 43899
rect 20329 43822 23210 43899
rect 20329 43758 22876 43822
rect 22940 43758 23210 43822
rect 20329 43701 23210 43758
rect 20130 43700 23210 43701
rect 25510 43612 25650 43670
rect 25510 43548 25558 43612
rect 25622 43548 25650 43612
rect 25510 43500 25650 43548
rect 20441 43340 20639 43345
rect 20440 43339 23850 43340
rect 20440 43141 20441 43339
rect 20639 43232 23850 43339
rect 20639 43168 23612 43232
rect 23676 43168 23850 43232
rect 20639 43141 23850 43168
rect 20440 43140 23850 43141
rect 20441 43135 20639 43140
rect 24348 42642 24412 42648
rect 25977 42640 26043 42643
rect 24412 42638 26043 42640
rect 24412 42582 25982 42638
rect 26038 42582 26043 42638
rect 24412 42580 26043 42582
rect 24348 42572 24412 42578
rect 25977 42577 26043 42580
rect 25078 42238 25084 42302
rect 25148 42300 25154 42302
rect 25757 42300 25823 42303
rect 25148 42298 25823 42300
rect 25148 42242 25762 42298
rect 25818 42242 25823 42298
rect 25148 42240 25823 42242
rect 25148 42238 25154 42240
rect 25757 42237 25823 42240
rect 25337 42020 25403 42023
rect 26556 42022 26620 42028
rect 25337 42018 26556 42020
rect 25337 41962 25342 42018
rect 25398 41962 26556 42018
rect 25337 41960 26556 41962
rect 25337 41957 25403 41960
rect 26556 41952 26620 41958
rect 25097 41840 25163 41843
rect 27292 41842 27356 41848
rect 25097 41838 27292 41840
rect 25097 41782 25102 41838
rect 25158 41782 27292 41838
rect 25097 41780 27292 41782
rect 25097 41777 25163 41780
rect 27292 41772 27356 41778
rect 24897 41660 24963 41663
rect 28028 41662 28092 41668
rect 19720 41630 19900 41660
rect 17684 41550 17690 41630
rect 17770 41550 19771 41630
rect 19851 41550 19900 41630
rect 24897 41658 28028 41660
rect 24897 41602 24902 41658
rect 24958 41602 28028 41658
rect 24897 41600 28028 41602
rect 24897 41597 24963 41600
rect 28028 41592 28092 41598
rect 19720 41530 19900 41550
rect 24697 41500 24763 41503
rect 28758 41500 28764 41502
rect 24697 41498 28764 41500
rect 24697 41442 24702 41498
rect 24758 41442 28764 41498
rect 24697 41440 28764 41442
rect 24697 41437 24763 41440
rect 28758 41438 28764 41440
rect 28828 41438 28834 41502
rect 19606 41380 19696 41385
rect 16970 41372 19611 41380
rect 16970 41308 16988 41372
rect 17052 41308 19611 41372
rect 16970 41300 19611 41308
rect 19691 41300 19696 41380
rect 24387 41370 24453 41373
rect 29500 41372 29564 41378
rect 24387 41368 29500 41370
rect 24387 41312 24392 41368
rect 24448 41312 29500 41368
rect 24387 41310 29500 41312
rect 24387 41307 24453 41310
rect 29500 41302 29564 41308
rect 19606 41295 19696 41300
rect 25375 28220 25985 28225
rect 16600 28215 25380 28220
rect 16600 27625 16605 28215
rect 17195 27625 25380 28215
rect 16600 27620 25380 27625
rect 25980 27620 25985 28220
rect 25375 27615 25985 27620
rect 28250 8938 31430 8970
rect 28250 8895 31050 8938
rect 28250 8785 28275 8895
rect 28385 8820 31050 8895
rect 31168 8900 31430 8938
rect 31168 8899 31432 8900
rect 31168 8820 31313 8899
rect 28385 8785 31313 8820
rect 28250 8781 31313 8785
rect 31431 8781 31437 8899
rect 28250 8780 31432 8781
rect 28250 8770 31430 8780
rect 28250 8760 31160 8770
rect 20410 7805 20670 7820
rect 20410 7595 20435 7805
rect 20645 7595 20670 7805
rect 20410 7580 20670 7595
rect 20110 7505 20350 7530
rect 20110 7295 20125 7505
rect 20335 7295 20350 7505
rect 20110 7280 20350 7295
rect 20235 1530 20545 1535
rect 20235 1230 20240 1530
rect 20540 1399 27340 1530
rect 20540 1281 26897 1399
rect 27015 1281 27340 1399
rect 20540 1230 27340 1281
rect 20235 1225 20545 1230
rect 19645 970 19955 975
rect 19645 670 19650 970
rect 19950 809 22810 970
rect 19950 691 22481 809
rect 22599 691 22810 809
rect 19950 670 22810 691
rect 19645 665 19955 670
<< via3 >>
rect 20131 43701 20329 43899
rect 22876 43758 22940 43822
rect 25558 43608 25622 43612
rect 25558 43552 25562 43608
rect 25562 43552 25618 43608
rect 25618 43552 25622 43608
rect 25558 43548 25622 43552
rect 20441 43141 20639 43339
rect 23612 43168 23676 43232
rect 24348 42578 24412 42642
rect 25084 42238 25148 42302
rect 26556 41958 26620 42022
rect 27292 41778 27356 41842
rect 17690 41550 17770 41630
rect 28028 41598 28092 41662
rect 28764 41438 28828 41502
rect 16988 41308 17052 41372
rect 29500 41308 29564 41372
rect 31050 8820 31168 8938
rect 31313 8781 31431 8899
rect 20435 7800 20645 7805
rect 20435 7600 20440 7800
rect 20440 7600 20640 7800
rect 20640 7600 20645 7800
rect 20435 7595 20645 7600
rect 20125 7500 20335 7505
rect 20125 7300 20130 7500
rect 20130 7300 20330 7500
rect 20330 7300 20335 7500
rect 20125 7295 20335 7300
rect 26897 1281 27015 1399
rect 22481 691 22599 809
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 200 1000 500 44152
rect 9800 1000 10100 44152
rect 16990 41373 17050 45152
rect 17726 42480 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 20130 43899 20330 43900
rect 20130 43701 20131 43899
rect 20329 43701 20330 43899
rect 22878 43823 22938 45152
rect 22875 43822 22941 43823
rect 22875 43758 22876 43822
rect 22940 43758 22941 43822
rect 22875 43757 22941 43758
rect 17690 42340 17830 42480
rect 17690 41631 17770 42340
rect 17689 41630 17771 41631
rect 17689 41550 17690 41630
rect 17770 41550 17771 41630
rect 17689 41549 17771 41550
rect 16987 41372 17053 41373
rect 16987 41308 16988 41372
rect 17052 41308 17053 41372
rect 16987 41307 17053 41308
rect 20130 7506 20330 43701
rect 20440 43339 20640 43340
rect 20440 43141 20441 43339
rect 20639 43141 20640 43339
rect 23614 43233 23674 45152
rect 23611 43232 23677 43233
rect 23611 43168 23612 43232
rect 23676 43168 23677 43232
rect 23611 43167 23677 43168
rect 20440 7806 20640 43141
rect 24350 42643 24410 45152
rect 24347 42642 24413 42643
rect 24347 42578 24348 42642
rect 24412 42578 24413 42642
rect 24347 42577 24413 42578
rect 25086 42303 25146 45152
rect 25557 43612 25623 43613
rect 25557 43548 25558 43612
rect 25622 43610 25623 43612
rect 25822 43610 25882 45152
rect 25622 43550 25882 43610
rect 25622 43548 25623 43550
rect 25557 43547 25623 43548
rect 25083 42302 25149 42303
rect 25083 42238 25084 42302
rect 25148 42238 25149 42302
rect 25083 42237 25149 42238
rect 26558 42023 26618 45152
rect 26555 42022 26621 42023
rect 26555 41958 26556 42022
rect 26620 41958 26621 42022
rect 26555 41957 26621 41958
rect 27294 41843 27354 45152
rect 27291 41842 27357 41843
rect 27291 41778 27292 41842
rect 27356 41778 27357 41842
rect 27291 41777 27357 41778
rect 28030 41663 28090 45152
rect 28027 41662 28093 41663
rect 28027 41598 28028 41662
rect 28092 41598 28093 41662
rect 28027 41597 28093 41598
rect 28766 41503 28826 45152
rect 28763 41502 28829 41503
rect 28763 41438 28764 41502
rect 28828 41438 28829 41502
rect 28763 41437 28829 41438
rect 29502 41373 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29499 41372 29565 41373
rect 29499 41308 29500 41372
rect 29564 41308 29565 41372
rect 29499 41307 29565 41308
rect 31050 8939 31430 8970
rect 31049 8938 31430 8939
rect 31049 8820 31050 8938
rect 31168 8900 31430 8938
rect 31168 8899 31432 8900
rect 31168 8820 31313 8899
rect 31049 8819 31313 8820
rect 31050 8781 31313 8819
rect 31431 8781 31432 8899
rect 20434 7805 20646 7806
rect 20434 7595 20435 7805
rect 20645 7595 20646 7805
rect 20434 7594 20646 7595
rect 20124 7505 20336 7506
rect 20124 7295 20125 7505
rect 20335 7295 20336 7505
rect 20124 7294 20336 7295
rect 26896 1399 27016 1400
rect 26896 1281 26897 1399
rect 27015 1281 27016 1399
rect 31050 1290 31432 8781
rect 22480 809 22600 810
rect 22480 691 22481 809
rect 22599 691 22600 809
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 691
rect 26896 0 27016 1281
rect 31300 280 31432 1290
rect 31312 0 31432 280
use gilbert_mixer  gilbert_mixer_0
timestamp 1716076243
transform 1 0 3010 0 1 31000
box -1010 -1000 6620 10400
use gilbert_mixer  gilbert_mixer_1
timestamp 1716076243
transform 1 0 22010 0 1 3000
box -1010 -1000 6620 10400
use idac1  idac1_0
timestamp 1717254928
transform 0 -1 25200 1 0 30638
box -1638 -3300 11376 3200
use pll1_dco  pll1_dco_0
timestamp 1717256045
transform 0 1 18771 -1 0 39032
box -2140 -740 2480 1250
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM2
timestamp 1713470961
transform 0 1 19139 -1 0 34676
box -296 -619 296 619
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
