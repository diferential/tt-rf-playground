magic
tech sky130A
magscale 1 2
timestamp 1713472767
<< nwell >>
rect -200 2630 990 2640
rect 360 1400 430 2630
<< pwell >>
rect 1140 2040 1800 2100
rect 1140 1380 1240 2040
rect 1680 1380 1800 2040
rect 1140 1300 1800 1380
rect 1140 1280 2000 1300
rect -400 1120 2000 1280
rect -400 480 -300 1120
rect 120 480 260 1120
rect 700 480 840 1120
rect 1280 480 1420 1120
rect 1840 480 2000 1120
rect -400 200 2000 480
<< psubdiff >>
rect 1700 1300 1800 2100
rect 1380 1220 1800 1240
rect -340 1140 1880 1220
rect 1380 1130 1880 1140
rect 1380 1120 1420 1130
rect 1830 1120 1880 1130
rect 1400 1090 1420 1120
<< locali >>
rect -400 2700 2000 2800
rect -400 1520 -340 2700
rect -220 2580 -180 2700
rect 940 2580 1060 2700
rect -220 2568 -68 2580
rect 260 2568 532 2580
rect 860 2568 1060 2580
rect -220 2540 1060 2568
rect -220 2506 -120 2540
rect -220 1532 -164 2506
rect -130 1532 -120 2506
rect -220 1520 -120 1532
rect -400 1480 -120 1520
rect 300 2506 480 2540
rect 300 1532 322 2506
rect 356 1532 436 2506
rect 470 1532 480 2506
rect 300 1480 480 1532
rect 900 2520 1060 2540
rect 1860 2520 2000 2700
rect 900 2506 2000 2520
rect 900 1532 922 2506
rect 956 2400 2000 2506
rect 956 1532 1020 2400
rect 900 1480 1020 1532
rect -400 1470 1020 1480
rect -400 1436 -68 1470
rect 260 1436 532 1470
rect 860 1436 1020 1470
rect -400 1420 1020 1436
rect 1140 2040 1800 2100
rect 1140 2020 1240 2040
rect 1140 1320 1160 2020
rect 1220 1380 1240 2020
rect 1680 2020 1800 2040
rect 1680 1380 1700 2020
rect 1220 1320 1700 1380
rect 1760 1320 1800 2020
rect 1140 1300 1800 1320
rect -400 1260 2000 1300
rect -400 1150 -340 1260
rect -400 1140 140 1150
rect 1860 1140 2000 1260
rect -400 1120 2000 1140
rect -400 1088 -300 1120
rect -400 532 -364 1088
rect -330 532 -300 1088
rect -400 480 -300 532
rect 120 1088 260 1120
rect 120 532 216 1088
rect 250 532 260 1088
rect 120 480 260 532
rect 700 480 840 1120
rect 1280 480 1420 1120
rect 1840 1088 2000 1120
rect 1840 532 1862 1088
rect 1896 532 2000 1088
rect 1840 480 2000 532
rect -400 440 2000 480
rect -400 300 -300 440
rect 1900 300 2000 440
rect -400 200 2000 300
<< viali >>
rect -340 1520 -220 2700
rect -180 2580 940 2700
rect -68 2568 260 2580
rect 532 2568 860 2580
rect -164 1532 -130 2506
rect 322 1532 356 2506
rect 436 1532 470 2506
rect 1060 2520 1860 2700
rect 922 1532 956 2506
rect -68 1436 260 1470
rect 532 1436 860 1470
rect 1160 1320 1220 2020
rect 1700 1320 1760 2020
rect -340 1150 1860 1260
rect 140 1140 1860 1150
rect -364 532 -330 1088
rect 216 532 250 1088
rect 1862 532 1896 1088
rect -300 300 1900 440
<< metal1 >>
rect -400 2700 2000 2800
rect -400 1520 -340 2700
rect -220 2580 -180 2700
rect 940 2580 1060 2700
rect -220 2568 -68 2580
rect 260 2568 532 2580
rect 860 2568 1060 2580
rect -220 2540 1060 2568
rect -220 2506 -120 2540
rect -220 1532 -164 2506
rect -130 1532 -120 2506
rect 220 2506 560 2540
rect 80 2480 140 2500
rect 40 2460 120 2480
rect -90 1660 -80 2020
rect 0 1660 10 2020
rect 60 1580 160 2460
rect 220 1620 322 2506
rect 40 1560 160 1580
rect 40 1540 140 1560
rect -220 1520 -120 1532
rect -400 1480 -120 1520
rect 240 1532 322 1620
rect 356 1532 436 2506
rect 470 1532 560 2506
rect 900 2520 1060 2540
rect 1860 2520 2000 2700
rect 900 2506 2000 2520
rect 640 2280 840 2500
rect 640 2220 680 2280
rect 760 2220 840 2280
rect 640 1540 840 2220
rect 240 1480 560 1532
rect 900 1532 922 2506
rect 956 2400 2000 2506
rect 956 1532 1020 2400
rect 900 1480 1020 1532
rect -400 1470 1020 1480
rect -400 1436 -68 1470
rect 260 1436 532 1470
rect 860 1436 1020 1470
rect -400 1420 1020 1436
rect 1140 2040 1800 2100
rect 1140 2020 1240 2040
rect 1140 1320 1160 2020
rect 1220 1380 1240 2020
rect 1680 2020 1800 2040
rect 1680 1380 1700 2020
rect 1220 1320 1700 1380
rect 1760 1320 1800 2020
rect 1140 1300 1800 1320
rect 1140 1280 2000 1300
rect -400 1260 2000 1280
rect -400 1150 -340 1260
rect -400 1140 140 1150
rect 1860 1140 2000 1260
rect -400 1088 -300 1140
rect 120 1120 2000 1140
rect -400 532 -364 1088
rect -330 532 -300 1088
rect -198 1048 -188 1100
rect -20 1048 -10 1100
rect 120 1088 260 1120
rect -400 480 -300 532
rect 120 532 216 1088
rect 250 532 260 1088
rect 120 480 260 532
rect 700 480 840 1120
rect 1280 480 1420 1120
rect 1840 1088 2000 1120
rect 1840 532 1862 1088
rect 1896 532 2000 1088
rect 1840 480 2000 532
rect -400 440 2000 480
rect -400 300 -300 440
rect 1900 300 2000 440
rect -400 200 2000 300
<< via1 >>
rect -80 1660 0 2020
rect 680 2220 760 2280
rect -188 1048 -20 1100
<< metal2 >>
rect -400 2300 -200 2360
rect 1800 2300 2000 2360
rect -400 2200 160 2300
rect 640 2280 2000 2300
rect 640 2220 680 2280
rect 760 2220 2000 2280
rect 640 2200 2000 2220
rect -400 2160 -200 2200
rect 1800 2160 2000 2200
rect -160 2020 80 2100
rect -160 1660 -80 2020
rect 0 1660 80 2020
rect -160 1260 80 1660
rect -240 1100 80 1260
rect -240 1048 -188 1100
rect -20 1048 80 1100
rect -240 980 80 1048
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM1
timestamp 1713470961
transform 1 0 96 0 1 2019
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM2
timestamp 1713470961
transform 1 0 696 0 1 2019
box -296 -619 296 619
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM3
timestamp 1713470961
transform 1 0 -104 0 1 810
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM4
timestamp 1713470961
transform 1 0 476 0 1 810
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM5
timestamp 1713470961
transform 1 0 1056 0 1 810
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM6
timestamp 1713470961
transform 1 0 1636 0 1 810
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM7
timestamp 1713470961
transform 1 0 1456 0 1 1700
box -296 -410 296 410
<< labels >>
flabel metal1 -400 2700 -300 2800 0 FreeSans 1600 0 0 0 VDD
port 5 nsew
<< end >>
