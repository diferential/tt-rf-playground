magic
tech sky130A
magscale 1 2
timestamp 1723341833
<< metal1 >>
rect 0 1160 660 1540
rect 1060 1360 2820 1540
rect 1400 1220 1480 1360
rect 2140 1220 2220 1360
rect 280 980 360 1160
rect 1260 1120 1740 1160
rect 1300 1020 1580 1060
rect 140 880 540 920
rect 1540 880 1580 1020
rect 180 800 460 840
rect 220 640 260 800
rect 0 580 260 640
rect 220 480 260 580
rect 500 620 540 880
rect 1530 820 1540 880
rect 1600 820 1610 880
rect 1540 780 1580 820
rect 1700 780 1740 1120
rect 1820 1120 2380 1160
rect 1820 880 1860 1120
rect 2040 1020 2320 1060
rect 2040 880 2080 1020
rect 1810 820 1820 880
rect 1880 820 1890 880
rect 2020 820 2080 880
rect 1540 720 1600 780
rect 1670 720 1680 780
rect 1740 720 1750 780
rect 500 580 1540 620
rect 210 420 220 480
rect 280 420 290 480
rect 220 380 260 420
rect 500 340 540 580
rect 1530 560 1540 580
rect 1600 560 1610 620
rect 590 440 600 500
rect 660 480 670 500
rect 660 440 1560 480
rect 1700 380 1740 720
rect 1100 340 1740 380
rect 1820 380 1860 820
rect 2040 780 2080 820
rect 2010 720 2020 780
rect 2080 720 2090 780
rect 2010 560 2020 620
rect 2080 560 2090 620
rect 2040 480 2080 560
rect 2000 440 2580 480
rect 1820 340 2480 380
rect 320 300 540 340
rect 140 100 220 300
rect 940 140 1600 240
rect 1960 140 2620 240
rect 780 100 2820 140
rect 0 0 2820 100
<< via1 >>
rect 1540 820 1600 880
rect 1820 820 1880 880
rect 1680 720 1740 780
rect 220 420 280 480
rect 1540 560 1600 620
rect 600 440 660 500
rect 2020 720 2080 780
rect 2020 560 2080 620
<< metal2 >>
rect 1540 880 1600 890
rect 1820 880 1880 890
rect 1600 820 1820 860
rect 2640 860 2740 920
rect 1880 820 2740 860
rect 1540 810 1600 820
rect 1820 810 1880 820
rect 1680 780 1740 790
rect 2020 780 2080 790
rect 1740 720 2020 760
rect 2080 720 2740 760
rect 1680 710 1740 720
rect 2020 710 2080 720
rect 2640 660 2740 720
rect 1540 620 1600 630
rect 2020 620 2080 630
rect 1600 580 2020 620
rect 1540 550 1600 560
rect 2020 550 2080 560
rect 600 500 660 510
rect 220 480 280 490
rect 280 440 600 480
rect 600 430 660 440
rect 220 410 280 420
use sky130_fd_pr__nfet_01v8_FETKPT  sky130_fd_pr__nfet_01v8_FETKPT_0
timestamp 1723339032
transform 1 0 266 0 1 279
box -246 -279 246 279
use sky130_fd_pr__nfet_01v8_PL5MMV  sky130_fd_pr__nfet_01v8_PL5MMV_0
timestamp 1723338882
transform 1 0 246 0 1 279
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_8MENFK  sky130_fd_pr__nfet_g5v0d10v5_8MENFK_0
timestamp 1723341670
transform 1 0 2295 0 1 327
box -515 -327 515 327
use sky130_fd_pr__nfet_g5v0d10v5_8MENFK  sky130_fd_pr__nfet_g5v0d10v5_8MENFK_1
timestamp 1723341670
transform 1 0 1275 0 1 327
box -515 -327 515 327
use sky130_fd_pr__pfet_01v8_lvt_3K87YT  sky130_fd_pr__pfet_01v8_lvt_3K87YT_0
timestamp 1723341670
transform 1 0 325 0 1 944
box -325 -284 325 284
use sky130_fd_pr__pfet_g5v0d10v5_3JABYW  sky130_fd_pr__pfet_g5v0d10v5_3JABYW_0
timestamp 1723341670
transform 1 0 2187 0 1 1182
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_3JABYW  sky130_fd_pr__pfet_g5v0d10v5_3JABYW_1
timestamp 1723341670
transform 1 0 1447 0 1 1182
box -387 -362 387 362
<< labels >>
flabel metal1 0 580 60 640 0 FreeSans 1600 0 0 0 D
port 1 nsew
flabel metal1 500 580 540 620 0 FreeSans 320 0 0 0 DB
flabel metal1 0 1160 80 1240 0 FreeSans 1600 0 0 0 VDDL
port 2 nsew
flabel metal1 0 0 80 80 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal1 2660 1360 2820 1540 0 FreeSans 1600 0 0 0 VDDH
port 5 nsew
flabel space 2640 820 2740 920 0 FreeSans 800 0 0 0 Q
port 7 nsew
flabel space 2640 660 2740 760 0 FreeSans 800 0 0 0 QB
port 8 nsew
<< end >>
