magic
tech sky130A
magscale 1 2
timestamp 1713067979
<< pwell >>
rect -683 -979 683 979
<< nmos >>
rect -487 -769 -287 831
rect -229 -769 -29 831
rect 29 -769 229 831
rect 287 -769 487 831
<< ndiff >>
rect -545 819 -487 831
rect -545 -757 -533 819
rect -499 -757 -487 819
rect -545 -769 -487 -757
rect -287 819 -229 831
rect -287 -757 -275 819
rect -241 -757 -229 819
rect -287 -769 -229 -757
rect -29 819 29 831
rect -29 -757 -17 819
rect 17 -757 29 819
rect -29 -769 29 -757
rect 229 819 287 831
rect 229 -757 241 819
rect 275 -757 287 819
rect 229 -769 287 -757
rect 487 819 545 831
rect 487 -757 499 819
rect 533 -757 545 819
rect 487 -769 545 -757
<< ndiffc >>
rect -533 -757 -499 819
rect -275 -757 -241 819
rect -17 -757 17 819
rect 241 -757 275 819
rect 499 -757 533 819
<< psubdiff >>
rect -647 909 647 943
rect -647 847 -613 909
rect 613 847 647 909
rect -647 -909 -613 -847
rect 613 -909 647 -847
rect -647 -943 -551 -909
rect 551 -943 647 -909
<< psubdiffcont >>
rect -647 -847 -613 847
rect 613 -847 647 847
rect -551 -943 551 -909
<< poly >>
rect -487 831 -287 857
rect -229 831 -29 857
rect 29 831 229 857
rect 287 831 487 857
rect -487 -807 -287 -769
rect -487 -841 -471 -807
rect -303 -841 -287 -807
rect -487 -857 -287 -841
rect -229 -807 -29 -769
rect -229 -841 -213 -807
rect -45 -841 -29 -807
rect -229 -857 -29 -841
rect 29 -807 229 -769
rect 29 -841 45 -807
rect 213 -841 229 -807
rect 29 -857 229 -841
rect 287 -807 487 -769
rect 287 -841 303 -807
rect 471 -841 487 -807
rect 287 -857 487 -841
<< polycont >>
rect -471 -841 -303 -807
rect -213 -841 -45 -807
rect 45 -841 213 -807
rect 303 -841 471 -807
<< locali >>
rect -647 847 -613 943
rect 613 847 647 943
rect -533 819 -499 835
rect -533 -773 -499 -757
rect -275 819 -241 835
rect -275 -773 -241 -757
rect -17 819 17 835
rect -17 -773 17 -757
rect 241 819 275 835
rect 241 -773 275 -757
rect 499 819 533 835
rect 499 -773 533 -757
rect -487 -841 -471 -807
rect -303 -841 -287 -807
rect -229 -841 -213 -807
rect -45 -841 -29 -807
rect 29 -841 45 -807
rect 213 -841 229 -807
rect 287 -841 303 -807
rect 471 -841 487 -807
rect -647 -943 -551 -909
rect 551 -943 647 -909
<< viali >>
rect -613 909 613 943
rect -647 -847 -613 -182
rect -533 172 -499 802
rect -275 -740 -241 -110
rect -17 172 17 802
rect 241 -740 275 -110
rect 499 172 533 802
rect -471 -841 -303 -807
rect -213 -841 -45 -807
rect 45 -841 213 -807
rect 303 -841 471 -807
rect -647 -909 -613 -847
rect 613 -847 647 -182
rect 613 -909 647 -847
<< metal1 >>
rect -625 943 625 949
rect -625 909 -613 943
rect 613 909 625 943
rect -625 903 625 909
rect -539 802 -493 814
rect -539 172 -533 802
rect -499 172 -493 802
rect -539 160 -493 172
rect -23 802 23 814
rect -23 172 -17 802
rect 17 172 23 802
rect -23 160 23 172
rect 493 802 539 814
rect 493 172 499 802
rect 533 172 539 802
rect 493 160 539 172
rect -281 -110 -235 -98
rect -653 -182 -607 -170
rect -653 -909 -647 -182
rect -613 -909 -607 -182
rect -281 -740 -275 -110
rect -241 -740 -235 -110
rect -281 -752 -235 -740
rect 235 -110 281 -98
rect 235 -740 241 -110
rect 275 -740 281 -110
rect 235 -752 281 -740
rect 607 -182 653 -170
rect -483 -807 -291 -801
rect -483 -841 -471 -807
rect -303 -841 -291 -807
rect -483 -847 -291 -841
rect -225 -807 -33 -801
rect -225 -841 -213 -807
rect -45 -841 -33 -807
rect -225 -847 -33 -841
rect 33 -807 225 -801
rect 33 -841 45 -807
rect 213 -841 225 -807
rect 33 -847 225 -841
rect 291 -807 483 -801
rect 291 -841 303 -807
rect 471 -841 483 -807
rect 291 -847 483 -841
rect -653 -921 -607 -909
rect 607 -909 613 -182
rect 647 -909 653 -182
rect 607 -921 653 -909
<< properties >>
string FIXED_BBOX -630 -926 630 926
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
