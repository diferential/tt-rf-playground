magic
tech sky130A
magscale 1 2
timestamp 1717271345
<< checkpaint >>
rect -3732 -3932 35702 49084
<< locali >>
rect 26650 30325 26950 30350
rect 26650 30075 26675 30325
rect 26925 30075 26950 30325
rect 26650 30050 26950 30075
rect 22400 25240 22560 26420
rect 22620 25990 22840 26300
rect 22620 25956 22683 25990
rect 22717 25956 22840 25990
rect 22620 25918 22840 25956
rect 22620 25884 22683 25918
rect 22717 25884 22840 25918
rect 22620 25846 22840 25884
rect 22620 25812 22683 25846
rect 22717 25812 22840 25846
rect 22620 25774 22840 25812
rect 22620 25740 22683 25774
rect 22717 25740 22840 25774
rect 22620 25330 22840 25740
<< viali >>
rect 26675 30075 26925 30325
rect 22683 25956 22717 25990
rect 22683 25884 22717 25918
rect 22683 25812 22717 25846
rect 22683 25740 22717 25774
<< metal1 >>
rect 19720 41616 19900 41660
rect 19720 41564 19785 41616
rect 19837 41564 19900 41616
rect 19720 41530 19900 41564
rect 19611 41366 19691 41386
rect 19611 41314 19625 41366
rect 19677 41314 19691 41366
rect 19211 41122 19411 41138
rect 16600 41110 16740 41116
rect 16600 41098 18171 41110
rect 16600 40982 16612 41098
rect 16728 40982 18171 41098
rect 16600 40970 18171 40982
rect 16600 40964 16740 40970
rect 18891 40938 19031 40950
rect 18891 40822 18903 40938
rect 19019 40822 19031 40938
rect 19211 40942 19221 41122
rect 19401 40942 19411 41122
rect 19611 41000 19691 41314
rect 19771 41000 19851 41530
rect 19211 40926 19411 40942
rect 18891 40810 19031 40822
rect 26600 30325 27000 30500
rect 22090 30290 22310 30300
rect 22090 30110 22110 30290
rect 22290 30110 22310 30290
rect 22090 30100 22310 30110
rect 26600 30075 26675 30325
rect 26925 30075 27000 30325
rect 26600 30000 27000 30075
rect 22390 29890 22610 29900
rect 22390 29710 22410 29890
rect 22590 29710 22610 29890
rect 22390 29700 22610 29710
rect 22090 29490 22310 29500
rect 22090 29310 22110 29490
rect 22290 29310 22310 29490
rect 22090 29300 22310 29310
rect 22400 25930 22560 26020
rect 22224 25908 22560 25930
rect 22224 25792 22252 25908
rect 22368 25792 22560 25908
rect 22224 25770 22560 25792
rect 22400 25740 22560 25770
rect 22620 25990 22850 26270
rect 22620 25956 22683 25990
rect 22717 25977 22850 25990
rect 22620 25925 22689 25956
rect 22741 25925 22850 25977
rect 22620 25918 22850 25925
rect 22620 25884 22683 25918
rect 22717 25913 22850 25918
rect 22620 25861 22689 25884
rect 22741 25861 22850 25913
rect 22620 25849 22850 25861
rect 22620 25846 22689 25849
rect 22620 25812 22683 25846
rect 22620 25797 22689 25812
rect 22741 25797 22850 25849
rect 22620 25785 22850 25797
rect 22620 25774 22689 25785
rect 22620 25740 22683 25774
rect 22620 25733 22689 25740
rect 22741 25733 22850 25785
rect 22620 25340 22850 25733
rect 21290 12872 21610 12900
rect 21290 12628 21328 12872
rect 21572 12628 21610 12872
rect 21290 12600 21610 12628
rect 22190 12872 22510 12900
rect 22190 12628 22228 12872
rect 22472 12628 22510 12872
rect 22190 12600 22510 12628
rect 21790 2390 22610 2400
rect 21790 2210 21822 2390
rect 22578 2210 22610 2390
rect 21790 2200 22610 2210
rect 24290 2372 24910 2400
rect 24290 2128 24318 2372
rect 24882 2128 24910 2372
rect 24290 2100 24910 2128
<< via1 >>
rect 19785 41564 19837 41616
rect 19625 41314 19677 41366
rect 16612 40982 16728 41098
rect 18903 40822 19019 40938
rect 19221 40942 19401 41122
rect 22110 30110 22290 30290
rect 26678 30078 26922 30322
rect 22410 29710 22590 29890
rect 22110 29310 22290 29490
rect 22252 25792 22368 25908
rect 22689 25956 22717 25977
rect 22717 25956 22741 25977
rect 22689 25925 22741 25956
rect 22689 25884 22717 25913
rect 22717 25884 22741 25913
rect 22689 25861 22741 25884
rect 22689 25846 22741 25849
rect 22689 25812 22717 25846
rect 22717 25812 22741 25846
rect 22689 25797 22741 25812
rect 22689 25774 22741 25785
rect 22689 25740 22717 25774
rect 22717 25740 22741 25774
rect 22689 25733 22741 25740
rect 21328 12628 21572 12872
rect 22228 12628 22472 12872
rect 21822 2210 22578 2390
rect 24318 2128 24882 2372
<< metal2 >>
rect 25530 43608 25630 43630
rect 25530 43552 25562 43608
rect 25618 43552 25630 43608
rect 25330 42018 25430 43170
rect 25330 41962 25342 42018
rect 25398 41962 25430 42018
rect 19720 41618 19900 41660
rect 19720 41562 19783 41618
rect 19839 41562 19900 41618
rect 19720 41530 19900 41562
rect 19590 41368 19710 41420
rect 19590 41312 19623 41368
rect 19679 41312 19710 41368
rect 19590 41290 19710 41312
rect 24390 41368 24450 41640
rect 24700 41498 24760 41690
rect 24900 41658 24960 41840
rect 25100 41838 25160 41950
rect 25330 41890 25430 41962
rect 25100 41782 25102 41838
rect 25158 41782 25160 41838
rect 25530 41830 25630 43552
rect 25730 42298 25830 43160
rect 25730 42242 25762 42298
rect 25818 42242 25830 42298
rect 25730 41900 25830 42242
rect 25950 42638 26050 43150
rect 25950 42582 25982 42638
rect 26038 42582 26050 42638
rect 25950 41914 26050 42582
rect 25100 41780 25160 41782
rect 25102 41773 25158 41780
rect 24900 41602 24902 41658
rect 24958 41602 24960 41658
rect 24900 41600 24960 41602
rect 24902 41593 24958 41600
rect 24693 41442 24702 41498
rect 24758 41442 24767 41498
rect 24700 41440 24760 41442
rect 24390 41312 24392 41368
rect 24448 41312 24450 41368
rect 24390 41310 24450 41312
rect 24392 41303 24448 41310
rect 19205 41122 19417 41132
rect 16594 41098 16746 41110
rect 16594 40982 16612 41098
rect 16728 40982 16746 41098
rect 16594 40970 16746 40982
rect 16600 28215 17200 40970
rect 18860 40948 19060 41020
rect 18860 40812 18893 40948
rect 19029 40812 19060 40948
rect 19205 40942 19221 41122
rect 19401 40942 19417 41122
rect 19205 40932 19417 40942
rect 18860 40780 19060 40812
rect 19211 40700 19411 40932
rect 19202 40668 19420 40700
rect 19202 40532 19243 40668
rect 19379 40532 19420 40668
rect 19202 40500 19420 40532
rect 26600 30322 27000 30500
rect 22100 30290 22300 30310
rect 22100 30110 22110 30290
rect 22290 30110 22300 30290
rect 22100 30090 22300 30110
rect 26600 30078 26678 30322
rect 26922 30078 27000 30322
rect 26600 30000 27000 30078
rect 22400 29890 22600 29910
rect 22400 29800 22410 29890
rect 22200 29710 22410 29800
rect 22590 29710 22600 29890
rect 22200 29690 22600 29710
rect 22200 29510 22400 29690
rect 22100 29490 22400 29510
rect 22100 29310 22110 29490
rect 22290 29310 22400 29490
rect 22100 29290 22400 29310
rect 16596 28188 17204 28215
rect 16596 27652 16632 28188
rect 17168 27652 17204 28188
rect 16596 27625 17204 27652
rect 16600 27620 17200 27625
rect 22200 26600 22400 29290
rect 23000 29000 23400 29800
rect 23000 26695 23200 29000
rect 25380 28188 25980 29838
rect 25380 27652 25412 28188
rect 25948 27652 25980 28188
rect 25380 27611 25980 27652
rect 22230 25908 22390 26600
rect 22230 25792 22252 25908
rect 22368 25792 22390 25908
rect 22230 25764 22390 25792
rect 22660 26585 23205 26695
rect 22660 25977 22770 26585
rect 22660 25925 22689 25977
rect 22741 25925 22770 25977
rect 22660 25913 22770 25925
rect 22660 25861 22689 25913
rect 22741 25861 22770 25913
rect 22660 25849 22770 25861
rect 22660 25797 22689 25849
rect 22741 25797 22770 25849
rect 22660 25785 22770 25797
rect 22660 25733 22689 25785
rect 22741 25733 22770 25785
rect 22660 24118 22770 25733
rect 22660 24062 22687 24118
rect 22743 24062 22770 24118
rect 22660 23960 22770 24062
rect 21300 12898 21600 12910
rect 21300 12602 21302 12898
rect 21598 12602 21600 12898
rect 21300 12590 21600 12602
rect 22200 12898 22500 12910
rect 22200 12602 22202 12898
rect 22498 12602 22500 12898
rect 22200 12590 22500 12602
rect 28275 8868 28385 8904
rect 28275 8812 28302 8868
rect 28358 8812 28385 8868
rect 28275 8776 28385 8812
rect 20431 7768 21230 7800
rect 20431 7632 20472 7768
rect 20608 7632 21230 7768
rect 20431 7600 21230 7632
rect 19990 7468 21220 7500
rect 19990 7332 20162 7468
rect 20298 7332 21220 7468
rect 19990 7300 21220 7332
rect 19650 4300 21320 4600
rect 19650 1000 19950 4300
rect 20240 3700 21310 4000
rect 20240 1528 20540 3700
rect 21800 2390 22600 2410
rect 21800 2368 21822 2390
rect 22578 2368 22600 2390
rect 21800 2232 21812 2368
rect 22588 2232 22600 2368
rect 21800 2210 21822 2232
rect 22578 2210 22600 2232
rect 21800 2190 22600 2210
rect 24300 2398 24900 2410
rect 24300 2372 24332 2398
rect 24868 2372 24900 2398
rect 24300 2128 24318 2372
rect 24882 2128 24900 2372
rect 24300 2102 24332 2128
rect 24868 2102 24900 2128
rect 24300 2090 24900 2102
rect 20240 1232 20242 1528
rect 20538 1232 20540 1528
rect 20240 1221 20540 1232
rect 19530 968 20000 1000
rect 19530 672 19652 968
rect 19948 672 20000 968
rect 19530 620 20000 672
<< via2 >>
rect 25562 43552 25618 43608
rect 25342 41962 25398 42018
rect 19783 41616 19839 41618
rect 19783 41564 19785 41616
rect 19785 41564 19837 41616
rect 19837 41564 19839 41616
rect 19783 41562 19839 41564
rect 19623 41366 19679 41368
rect 19623 41314 19625 41366
rect 19625 41314 19677 41366
rect 19677 41314 19679 41366
rect 19623 41312 19679 41314
rect 25102 41782 25158 41838
rect 25762 42242 25818 42298
rect 25982 42582 26038 42638
rect 24902 41602 24958 41658
rect 24702 41442 24758 41498
rect 24392 41312 24448 41368
rect 18893 40938 19029 40948
rect 18893 40822 18903 40938
rect 18903 40822 19019 40938
rect 19019 40822 19029 40938
rect 18893 40812 19029 40822
rect 19243 40532 19379 40668
rect 22132 30132 22268 30268
rect 26692 30092 26908 30308
rect 22432 29732 22568 29868
rect 22132 29332 22268 29468
rect 16632 27652 17168 28188
rect 25412 27652 25948 28188
rect 22687 24062 22743 24118
rect 21302 12872 21598 12898
rect 21302 12628 21328 12872
rect 21328 12628 21572 12872
rect 21572 12628 21598 12872
rect 21302 12602 21598 12628
rect 22202 12872 22498 12898
rect 22202 12628 22228 12872
rect 22228 12628 22472 12872
rect 22472 12628 22498 12872
rect 22202 12602 22498 12628
rect 28302 8812 28358 8868
rect 20472 7632 20608 7768
rect 20162 7332 20298 7468
rect 21812 2232 21822 2368
rect 21822 2232 22578 2368
rect 22578 2232 22588 2368
rect 24332 2372 24868 2398
rect 24332 2128 24868 2372
rect 24332 2102 24868 2128
rect 20242 1232 20538 1528
rect 19652 672 19948 968
<< metal3 >>
rect 9331 44152 9629 44157
rect 710 44114 9630 44152
rect 10371 44150 10669 44155
rect 710 44032 9368 44114
rect 710 44012 2268 44032
rect 710 43948 796 44012
rect 860 43948 1532 44012
rect 1596 43968 2268 44012
rect 2332 43968 3004 44032
rect 3068 44012 4476 44032
rect 3068 43968 3740 44012
rect 1596 43948 3740 43968
rect 3804 43968 4476 44012
rect 4540 43968 5212 44032
rect 5276 43968 5948 44032
rect 6012 44012 9368 44032
rect 6012 43968 6688 44012
rect 3804 43948 6688 43968
rect 6752 43948 9368 44012
rect 710 43890 9368 43948
rect 9592 43890 9630 44114
rect 710 43852 9630 43890
rect 10370 44146 16430 44150
rect 16490 44146 16690 44150
rect 10370 44112 16690 44146
rect 10370 43888 10408 44112
rect 10632 44032 16690 44112
rect 10632 43968 12572 44032
rect 12636 43968 13308 44032
rect 13372 43968 14044 44032
rect 14108 43968 14780 44032
rect 14844 43968 15516 44032
rect 15580 44012 16690 44032
rect 15580 43968 16252 44012
rect 10632 43948 16252 43968
rect 16316 43948 16690 44012
rect 10632 43888 16690 43948
rect 20130 43899 23210 43900
rect 9331 43847 9629 43852
rect 10370 43850 16690 43888
rect 20125 43872 23210 43899
rect 10371 43845 10669 43850
rect 16320 43832 16520 43850
rect 20125 43728 20158 43872
rect 20302 43822 23210 43872
rect 20302 43758 22876 43822
rect 22940 43758 23210 43822
rect 20302 43728 23210 43758
rect 20125 43701 23210 43728
rect 20130 43700 23210 43701
rect 25510 43612 25650 43670
rect 25510 43548 25558 43612
rect 25622 43548 25650 43612
rect 25510 43500 25650 43548
rect 20441 43340 20639 43345
rect 20440 43312 23850 43340
rect 20440 43168 20468 43312
rect 20612 43232 23850 43312
rect 20612 43168 23612 43232
rect 23676 43168 23850 43232
rect 20440 43140 23850 43168
rect 20441 43135 20639 43140
rect 24348 42642 24412 42648
rect 25977 42640 26043 42643
rect 24412 42638 26043 42640
rect 24412 42582 25982 42638
rect 26038 42582 26043 42638
rect 24412 42580 26043 42582
rect 24348 42572 24412 42578
rect 25977 42577 26043 42580
rect 25078 42238 25084 42302
rect 25148 42300 25154 42302
rect 25757 42300 25823 42303
rect 25148 42298 25823 42300
rect 25148 42242 25762 42298
rect 25818 42242 25823 42298
rect 25148 42240 25823 42242
rect 25148 42238 25154 42240
rect 25757 42237 25823 42240
rect 25337 42020 25403 42023
rect 26556 42022 26620 42028
rect 25337 42018 26556 42020
rect 25337 41962 25342 42018
rect 25398 41962 26556 42018
rect 25337 41960 26556 41962
rect 25337 41957 25403 41960
rect 26556 41952 26620 41958
rect 25097 41840 25163 41843
rect 27292 41842 27356 41848
rect 25097 41838 27292 41840
rect 25097 41782 25102 41838
rect 25158 41782 27292 41838
rect 25097 41780 27292 41782
rect 25097 41777 25163 41780
rect 27292 41772 27356 41778
rect 24897 41660 24963 41663
rect 28028 41662 28092 41668
rect 19720 41630 19900 41660
rect 17684 41622 19900 41630
rect 17684 41558 17698 41622
rect 17762 41618 19900 41622
rect 17762 41562 19783 41618
rect 19839 41562 19900 41618
rect 24897 41658 28028 41660
rect 24897 41602 24902 41658
rect 24958 41602 28028 41658
rect 24897 41600 28028 41602
rect 24897 41597 24963 41600
rect 28028 41592 28092 41598
rect 17762 41558 19900 41562
rect 17684 41550 19900 41558
rect 19720 41530 19900 41550
rect 24697 41500 24763 41503
rect 28758 41500 28764 41502
rect 24697 41498 28764 41500
rect 24697 41442 24702 41498
rect 24758 41442 28764 41498
rect 24697 41440 28764 41442
rect 24697 41437 24763 41440
rect 28758 41438 28764 41440
rect 28828 41438 28834 41502
rect 19606 41380 19696 41385
rect 16970 41372 19696 41380
rect 16970 41308 16988 41372
rect 17052 41368 19696 41372
rect 17052 41312 19623 41368
rect 19679 41312 19696 41368
rect 17052 41308 19696 41312
rect 16970 41300 19696 41308
rect 24387 41370 24453 41373
rect 29500 41372 29564 41378
rect 24387 41368 29500 41370
rect 24387 41312 24392 41368
rect 24448 41312 29500 41368
rect 24387 41310 29500 41312
rect 24387 41307 24453 41310
rect 29500 41302 29564 41308
rect 19606 41295 19696 41300
rect 820 40972 1520 41100
rect 820 40908 928 40972
rect 992 40908 1008 40972
rect 1072 40950 1520 40972
rect 18886 40950 19036 40955
rect 1072 40948 19036 40950
rect 1072 40908 18893 40948
rect 820 40892 18893 40908
rect 820 40828 1228 40892
rect 1292 40828 1308 40892
rect 1372 40828 18893 40892
rect 820 40812 18893 40828
rect 19029 40812 19036 40948
rect 820 40810 19036 40812
rect 820 40632 1520 40810
rect 18886 40805 19036 40810
rect 19206 40700 19416 40705
rect 820 40568 1188 40632
rect 1252 40568 1268 40632
rect 1332 40568 1520 40632
rect 820 40460 1520 40568
rect 10794 40672 19416 40700
rect 10794 40528 10828 40672
rect 10972 40668 19416 40672
rect 10972 40532 19243 40668
rect 19379 40532 19416 40668
rect 10972 40528 19416 40532
rect 10794 40500 19416 40528
rect 19206 40495 19416 40500
rect 10551 32050 10849 32055
rect 10500 32012 21456 32050
rect 10500 31788 10588 32012
rect 10812 31788 21188 32012
rect 21412 31788 21456 32012
rect 10500 31750 21456 31788
rect 10551 31745 10849 31750
rect 22000 30268 22800 30400
rect 22000 30132 22132 30268
rect 22268 30132 22800 30268
rect 22000 29868 22800 30132
rect 26600 30312 27000 30500
rect 26600 30088 26688 30312
rect 26912 30088 27000 30312
rect 26600 30000 27000 30088
rect 22000 29732 22432 29868
rect 22568 29732 22800 29868
rect 951 29550 1249 29555
rect 22000 29550 22800 29732
rect 950 29512 22800 29550
rect 950 29288 988 29512
rect 1212 29468 22800 29512
rect 1212 29332 22132 29468
rect 22268 29332 22800 29468
rect 1212 29288 22800 29332
rect 950 29250 22800 29288
rect 951 29245 1249 29250
rect 22000 29200 22800 29250
rect 25375 28220 25985 28225
rect 16600 28188 25985 28220
rect 16600 27652 16632 28188
rect 17168 27652 25412 28188
rect 25948 27652 25985 28188
rect 16600 27620 25985 27652
rect 25375 27615 25985 27620
rect 17940 24172 22840 24200
rect 17940 24028 18008 24172
rect 18152 24118 22840 24172
rect 18152 24062 22687 24118
rect 22743 24062 22840 24118
rect 18152 24028 22840 24062
rect 17940 24000 22840 24028
rect 21100 12898 23100 13300
rect 851 12850 1149 12855
rect 21100 12850 21302 12898
rect 850 12812 21302 12850
rect 850 12588 888 12812
rect 1112 12602 21302 12812
rect 21598 12602 22202 12898
rect 22498 12602 23100 12898
rect 1112 12588 23100 12602
rect 850 12550 23100 12588
rect 851 12545 1149 12550
rect 21100 12200 23100 12550
rect 28250 8911 31430 8970
rect 28250 8868 31077 8911
rect 28250 8812 28302 8868
rect 28358 8847 31077 8868
rect 31141 8900 31430 8911
rect 31141 8899 31432 8900
rect 31141 8872 31437 8899
rect 31141 8847 31340 8872
rect 28358 8812 31340 8847
rect 28250 8808 31340 8812
rect 31404 8808 31437 8872
rect 28250 8781 31437 8808
rect 28250 8780 31432 8781
rect 28250 8770 31430 8780
rect 28250 8760 31160 8770
rect 20410 7772 20670 7820
rect 20410 7628 20468 7772
rect 20612 7628 20670 7772
rect 20410 7580 20670 7628
rect 20110 7472 20350 7530
rect 20110 7328 20158 7472
rect 20302 7328 20350 7472
rect 20110 7280 20350 7328
rect 21010 2490 25400 2500
rect 10541 2420 10839 2425
rect 21010 2420 25460 2490
rect 10540 2398 25460 2420
rect 10540 2382 24332 2398
rect 10540 2158 10578 2382
rect 10802 2368 24332 2382
rect 10802 2232 21812 2368
rect 22588 2232 24332 2368
rect 10802 2158 24332 2232
rect 10540 2120 24332 2158
rect 10541 2115 10839 2120
rect 21010 2102 24332 2120
rect 24868 2102 25460 2398
rect 21010 2000 25460 2102
rect 23900 1950 25460 2000
rect 20235 1530 20545 1535
rect 20235 1528 27340 1530
rect 20235 1232 20242 1528
rect 20538 1372 27340 1528
rect 20538 1308 26924 1372
rect 26988 1308 27340 1372
rect 20538 1232 27340 1308
rect 20235 1230 27340 1232
rect 20235 1225 20545 1230
rect 19645 970 19955 975
rect 19645 968 22810 970
rect 19645 672 19652 968
rect 19948 782 22810 968
rect 19948 718 22508 782
rect 22572 718 22810 782
rect 19948 672 22810 718
rect 19645 670 22810 672
rect 19645 665 19955 670
<< via3 >>
rect 796 43948 860 44012
rect 1532 43948 1596 44012
rect 2268 43968 2332 44032
rect 3004 43968 3068 44032
rect 3740 43948 3804 44012
rect 4476 43968 4540 44032
rect 5212 43968 5276 44032
rect 5948 43968 6012 44032
rect 6688 43948 6752 44012
rect 9368 43890 9592 44114
rect 10408 43888 10632 44112
rect 12572 43968 12636 44032
rect 13308 43968 13372 44032
rect 14044 43968 14108 44032
rect 14780 43968 14844 44032
rect 15516 43968 15580 44032
rect 16252 43948 16316 44012
rect 20158 43728 20302 43872
rect 22876 43758 22940 43822
rect 25558 43608 25622 43612
rect 25558 43552 25562 43608
rect 25562 43552 25618 43608
rect 25618 43552 25622 43608
rect 25558 43548 25622 43552
rect 20468 43168 20612 43312
rect 23612 43168 23676 43232
rect 24348 42578 24412 42642
rect 25084 42238 25148 42302
rect 26556 41958 26620 42022
rect 27292 41778 27356 41842
rect 17698 41558 17762 41622
rect 28028 41598 28092 41662
rect 28764 41438 28828 41502
rect 16988 41308 17052 41372
rect 29500 41308 29564 41372
rect 928 40908 992 40972
rect 1008 40908 1072 40972
rect 1228 40828 1292 40892
rect 1308 40828 1372 40892
rect 1188 40568 1252 40632
rect 1268 40568 1332 40632
rect 10828 40528 10972 40672
rect 10588 31788 10812 32012
rect 21188 31788 21412 32012
rect 26688 30308 26912 30312
rect 26688 30092 26692 30308
rect 26692 30092 26908 30308
rect 26908 30092 26912 30308
rect 26688 30088 26912 30092
rect 988 29288 1212 29512
rect 18008 24028 18152 24172
rect 888 12588 1112 12812
rect 31077 8847 31141 8911
rect 31340 8808 31404 8872
rect 20468 7768 20612 7772
rect 20468 7632 20472 7768
rect 20472 7632 20608 7768
rect 20608 7632 20612 7768
rect 20468 7628 20612 7632
rect 20158 7468 20302 7472
rect 20158 7332 20162 7468
rect 20162 7332 20298 7468
rect 20298 7332 20302 7468
rect 20158 7328 20302 7332
rect 10578 2158 10802 2382
rect 26924 1308 26988 1372
rect 22508 718 22572 782
<< metal4 >>
rect 200 40970 500 44152
rect 798 44013 858 45152
rect 1534 44013 1594 45152
rect 2270 44033 2330 45152
rect 3006 44033 3066 45152
rect 2267 44032 2333 44033
rect 795 44012 861 44013
rect 795 43948 796 44012
rect 860 43948 861 44012
rect 795 43947 861 43948
rect 1531 44012 1597 44013
rect 1531 43948 1532 44012
rect 1596 43948 1597 44012
rect 2267 43968 2268 44032
rect 2332 43968 2333 44032
rect 2267 43967 2333 43968
rect 3003 44032 3069 44033
rect 3003 43968 3004 44032
rect 3068 43968 3069 44032
rect 3742 44013 3802 45152
rect 4478 44033 4538 45152
rect 5214 44033 5274 45152
rect 5950 44033 6010 45152
rect 6686 45012 6746 45152
rect 7422 45012 7482 45152
rect 8158 45012 8218 45152
rect 8894 45012 8954 45152
rect 9630 45012 9690 45152
rect 10366 45012 10426 45152
rect 11102 45012 11162 45152
rect 11838 45012 11898 45152
rect 6686 44952 11898 45012
rect 4475 44032 4541 44033
rect 3003 43967 3069 43968
rect 3739 44012 3805 44013
rect 1531 43947 1597 43948
rect 3739 43948 3740 44012
rect 3804 43948 3805 44012
rect 4475 43968 4476 44032
rect 4540 43968 4541 44032
rect 4475 43967 4541 43968
rect 5211 44032 5277 44033
rect 5211 43968 5212 44032
rect 5276 43968 5277 44032
rect 5211 43967 5277 43968
rect 5947 44032 6013 44033
rect 5947 43968 5948 44032
rect 6012 43968 6013 44032
rect 6690 44013 6750 44952
rect 9330 44150 10100 44152
rect 9330 44114 10670 44150
rect 5947 43967 6013 43968
rect 6687 44012 6753 44013
rect 3739 43947 3805 43948
rect 6687 43948 6688 44012
rect 6752 43948 6753 44012
rect 6687 43947 6753 43948
rect 9330 43890 9368 44114
rect 9592 44112 10670 44114
rect 9592 43890 10408 44112
rect 9330 43888 10408 43890
rect 10632 43888 10670 44112
rect 12574 44033 12634 45152
rect 13310 44033 13370 45152
rect 14046 44033 14106 45152
rect 14782 44033 14842 45152
rect 15518 44033 15578 45152
rect 12571 44032 12637 44033
rect 12571 43968 12572 44032
rect 12636 43968 12637 44032
rect 12571 43967 12637 43968
rect 13307 44032 13373 44033
rect 13307 43968 13308 44032
rect 13372 43968 13373 44032
rect 13307 43967 13373 43968
rect 14043 44032 14109 44033
rect 14043 43968 14044 44032
rect 14108 43968 14109 44032
rect 14043 43967 14109 43968
rect 14779 44032 14845 44033
rect 14779 43968 14780 44032
rect 14844 43968 14845 44032
rect 14779 43967 14845 43968
rect 15515 44032 15581 44033
rect 15515 43968 15516 44032
rect 15580 43968 15581 44032
rect 16254 44013 16314 45152
rect 15515 43967 15581 43968
rect 16251 44012 16317 44013
rect 16251 43948 16252 44012
rect 16316 43948 16317 44012
rect 16251 43947 16317 43948
rect 9330 43852 10670 43888
rect 9800 43850 10670 43852
rect 820 40972 1520 41100
rect 820 40970 928 40972
rect 200 40908 928 40970
rect 992 40908 1008 40972
rect 1072 40908 1520 40972
rect 200 40892 1520 40908
rect 200 40828 1228 40892
rect 1292 40828 1308 40892
rect 1372 40828 1520 40892
rect 200 40670 1520 40828
rect 200 29550 500 40670
rect 820 40632 1520 40670
rect 820 40568 1188 40632
rect 1252 40568 1268 40632
rect 1332 40568 1520 40632
rect 820 40460 1520 40568
rect 9800 40700 10100 43850
rect 16990 41373 17050 45152
rect 17726 42480 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 20130 43872 20330 43900
rect 20130 43728 20158 43872
rect 20302 43728 20330 43872
rect 22878 43823 22938 45152
rect 22875 43822 22941 43823
rect 22875 43758 22876 43822
rect 22940 43758 22941 43822
rect 22875 43757 22941 43758
rect 17690 42340 17830 42480
rect 17690 41631 17770 42340
rect 17689 41622 17771 41631
rect 17689 41558 17698 41622
rect 17762 41558 17771 41622
rect 17689 41549 17771 41558
rect 16987 41372 17053 41373
rect 16987 41308 16988 41372
rect 17052 41308 17053 41372
rect 16987 41307 17053 41308
rect 10799 40700 11001 40701
rect 9800 40672 11001 40700
rect 9800 40528 10828 40672
rect 10972 40528 11001 40672
rect 9800 40500 11001 40528
rect 9800 32050 10100 40500
rect 10799 40499 11001 40500
rect 9800 32012 10850 32050
rect 9800 31788 10588 32012
rect 10812 31788 10850 32012
rect 9800 31750 10850 31788
rect 200 29512 1250 29550
rect 200 29288 988 29512
rect 1212 29288 1250 29512
rect 200 29250 1250 29288
rect 200 12850 500 29250
rect 200 12812 1150 12850
rect 200 12588 888 12812
rect 1112 12588 1150 12812
rect 200 12550 1150 12588
rect 200 4206 500 12550
rect 2436 5718 5828 6018
rect 2436 4206 2736 5718
rect 200 3906 2736 4206
rect 3918 3962 4218 5718
rect 5528 3998 5828 5718
rect 200 1000 500 3906
rect 2436 3218 2736 3906
rect 2436 2918 5756 3218
rect 5456 2504 5756 2918
rect 3918 2204 5756 2504
rect 9800 2420 10100 31750
rect 17979 24172 18181 24201
rect 17979 24028 18008 24172
rect 18152 24028 18181 24172
rect 17979 23999 18181 24028
rect 9800 2382 10840 2420
rect 5400 1608 5700 2204
rect 2582 1308 5700 1608
rect 9800 2158 10578 2382
rect 10802 2158 10840 2382
rect 9800 2120 10840 2158
rect 2582 894 2882 1308
rect 9800 1000 10100 2120
rect 17980 1064 18180 23999
rect 20130 7506 20330 43728
rect 20440 43312 20640 43340
rect 20440 43168 20468 43312
rect 20612 43168 20640 43312
rect 23614 43233 23674 45152
rect 20440 7806 20640 43168
rect 23611 43232 23677 43233
rect 23611 43168 23612 43232
rect 23676 43168 23677 43232
rect 23611 43167 23677 43168
rect 24350 42643 24410 45152
rect 24347 42642 24413 42643
rect 24347 42578 24348 42642
rect 24412 42578 24413 42642
rect 24347 42577 24413 42578
rect 25086 42303 25146 45152
rect 25557 43612 25623 43613
rect 25557 43548 25558 43612
rect 25622 43610 25623 43612
rect 25822 43610 25882 45152
rect 25622 43550 25882 43610
rect 25622 43548 25623 43550
rect 25557 43547 25623 43548
rect 25083 42302 25149 42303
rect 25083 42238 25084 42302
rect 25148 42238 25149 42302
rect 25083 42237 25149 42238
rect 26558 42023 26618 45152
rect 26555 42022 26621 42023
rect 26555 41958 26556 42022
rect 26620 41958 26621 42022
rect 26555 41957 26621 41958
rect 27294 41843 27354 45152
rect 27291 41842 27357 41843
rect 27291 41778 27292 41842
rect 27356 41778 27357 41842
rect 27291 41777 27357 41778
rect 28030 41663 28090 45152
rect 28027 41662 28093 41663
rect 28027 41598 28028 41662
rect 28092 41598 28093 41662
rect 28027 41597 28093 41598
rect 28766 41503 28826 45152
rect 28763 41502 28829 41503
rect 28763 41438 28764 41502
rect 28828 41438 28829 41502
rect 28763 41437 28829 41438
rect 29502 41373 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29499 41372 29565 41373
rect 29499 41308 29500 41372
rect 29564 41308 29565 41372
rect 29499 41307 29565 41308
rect 21149 32050 21451 32051
rect 21149 32012 26950 32050
rect 21149 31788 21188 32012
rect 21412 31788 26950 32012
rect 21149 31750 26950 31788
rect 21149 31749 21451 31750
rect 26650 30500 26950 31750
rect 26600 30312 27000 30500
rect 26600 30088 26688 30312
rect 26912 30088 27000 30312
rect 26600 30000 27000 30088
rect 31050 8939 31430 8970
rect 31049 8911 31430 8939
rect 31049 8847 31077 8911
rect 31141 8900 31430 8911
rect 31141 8872 31432 8900
rect 31141 8847 31340 8872
rect 31049 8819 31340 8847
rect 31050 8808 31340 8819
rect 31404 8808 31432 8872
rect 20434 7772 20646 7806
rect 20434 7628 20468 7772
rect 20612 7628 20646 7772
rect 20434 7594 20646 7628
rect 20124 7472 20336 7506
rect 20124 7328 20158 7472
rect 20302 7328 20336 7472
rect 20124 7294 20336 7328
rect 26866 1372 27046 1446
rect 26866 1308 26924 1372
rect 26988 1308 27046 1372
rect 2582 594 5590 894
rect 17980 322 18214 1064
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 322
rect 22450 782 22630 828
rect 22450 718 22508 782
rect 22572 718 22630 782
rect 22450 0 22630 718
rect 26866 0 27046 1308
rect 31050 1290 31432 8808
rect 31300 678 31432 1290
rect 31282 0 31462 678
use gilbert_mixer  gilbert_mixer_1
timestamp 1716061843
transform 1 0 22010 0 1 3000
box -1010 -1000 6620 10400
use idac1  idac1_0
timestamp 1717240528
transform 0 -1 25200 1 0 30638
box -1638 -3300 11376 3200
use pll1_dco  pll1_dco_0
timestamp 1717241645
transform 0 1 18771 -1 0 39032
box -2140 -740 2480 1250
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM2
timestamp 1713456561
transform -1 0 22696 0 -1 25819
box -296 -619 296 619
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 600 90 0 0 clk
port 1 nsew
flabel metal4 s 31004 45052 31004 45052 0 FreeSans 600 90 0 0 clk
flabel metal4 s 31004 45052 31004 45052 0 FreeSans 600 90 0 0 clk
flabel metal4 s 31004 45052 31004 45052 0 FreeSans 600 90 0 0 clk
flabel metal4 s 31004 45052 31004 45052 0 FreeSans 600 90 0 0 clk
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 600 90 0 0 ena
port 2 nsew
flabel metal4 s 31740 45052 31740 45052 0 FreeSans 600 90 0 0 ena
flabel metal4 s 31740 45052 31740 45052 0 FreeSans 600 90 0 0 ena
flabel metal4 s 31740 45052 31740 45052 0 FreeSans 600 90 0 0 ena
flabel metal4 s 31740 45052 31740 45052 0 FreeSans 600 90 0 0 ena
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 600 90 0 0 rst_n
port 3 nsew
flabel metal4 s 30268 45052 30268 45052 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 30268 45052 30268 45052 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 30268 45052 30268 45052 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 30268 45052 30268 45052 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 31282 0 31462 200 0 FreeSans 1200 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26866 0 27046 200 0 FreeSans 1200 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 26956 100 26956 100 0 FreeSans 1200 0 0 0 ua[1]
flabel metal4 s 22450 0 22630 200 0 FreeSans 1200 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 22540 100 22540 100 0 FreeSans 1200 0 0 0 ua[2]
flabel metal4 s 18034 0 18214 200 0 FreeSans 1200 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 18124 100 18124 100 0 FreeSans 1200 0 0 0 ua[3]
flabel metal4 s 13618 0 13798 200 0 FreeSans 1200 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 13708 100 13708 100 0 FreeSans 1200 0 0 0 ua[4]
flabel metal4 s 9202 0 9382 200 0 FreeSans 1200 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 9292 100 9292 100 0 FreeSans 1200 0 0 0 ua[5]
flabel metal4 s 4786 0 4966 200 0 FreeSans 1200 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 4876 100 4876 100 0 FreeSans 1200 0 0 0 ua[6]
flabel metal4 s 370 0 550 200 0 FreeSans 1200 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 460 100 460 100 0 FreeSans 1200 0 0 0 ua[7]
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 600 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 29532 45052 29532 45052 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 29532 45052 29532 45052 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 29532 45052 29532 45052 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 29532 45052 29532 45052 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 28796 45052 28796 45052 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 28796 45052 28796 45052 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 28796 45052 28796 45052 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 28796 45052 28796 45052 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 600 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 28060 45052 28060 45052 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 28060 45052 28060 45052 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 28060 45052 28060 45052 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 28060 45052 28060 45052 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 600 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 27324 45052 27324 45052 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 27324 45052 27324 45052 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 27324 45052 27324 45052 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 27324 45052 27324 45052 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 26588 45052 26588 45052 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 26588 45052 26588 45052 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 26588 45052 26588 45052 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 26588 45052 26588 45052 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 600 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 25852 45052 25852 45052 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 25852 45052 25852 45052 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 25852 45052 25852 45052 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 25852 45052 25852 45052 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 600 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 25116 45052 25116 45052 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 25116 45052 25116 45052 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 25116 45052 25116 45052 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 25116 45052 25116 45052 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 24380 45052 24380 45052 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 24380 45052 24380 45052 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 24380 45052 24380 45052 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 24380 45052 24380 45052 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 600 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 23644 45052 23644 45052 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 23644 45052 23644 45052 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 23644 45052 23644 45052 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 23644 45052 23644 45052 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 600 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 22908 45052 22908 45052 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22908 45052 22908 45052 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22908 45052 22908 45052 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22908 45052 22908 45052 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 22172 45052 22172 45052 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 22172 45052 22172 45052 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 22172 45052 22172 45052 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 22172 45052 22172 45052 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 600 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 21436 45052 21436 45052 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 21436 45052 21436 45052 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 21436 45052 21436 45052 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 21436 45052 21436 45052 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 600 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 20700 45052 20700 45052 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 20700 45052 20700 45052 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 20700 45052 20700 45052 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 20700 45052 20700 45052 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 19964 45052 19964 45052 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 19964 45052 19964 45052 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 19964 45052 19964 45052 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 19964 45052 19964 45052 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 600 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 19228 45052 19228 45052 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 19228 45052 19228 45052 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 19228 45052 19228 45052 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 19228 45052 19228 45052 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 600 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 18492 45052 18492 45052 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 18492 45052 18492 45052 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 18492 45052 18492 45052 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 18492 45052 18492 45052 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 600 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 5980 45052 5980 45052 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 5980 45052 5980 45052 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 5980 45052 5980 45052 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 5980 45052 5980 45052 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 600 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 5244 45052 5244 45052 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 5244 45052 5244 45052 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 5244 45052 5244 45052 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 5244 45052 5244 45052 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 600 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 4508 45052 4508 45052 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 4508 45052 4508 45052 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 4508 45052 4508 45052 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 4508 45052 4508 45052 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 600 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 3772 45052 3772 45052 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 3772 45052 3772 45052 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 3772 45052 3772 45052 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 3772 45052 3772 45052 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 600 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 3036 45052 3036 45052 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 3036 45052 3036 45052 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 3036 45052 3036 45052 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 3036 45052 3036 45052 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 600 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 2300 45052 2300 45052 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 2300 45052 2300 45052 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 2300 45052 2300 45052 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 2300 45052 2300 45052 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 600 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 1564 45052 1564 45052 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 1564 45052 1564 45052 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 1564 45052 1564 45052 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 1564 45052 1564 45052 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 798 44952 858 45152 0 FreeSans 600 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 828 45052 828 45052 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 828 45052 828 45052 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 828 45052 828 45052 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 828 45052 828 45052 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 600 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 11868 45052 11868 45052 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 11868 45052 11868 45052 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 11868 45052 11868 45052 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 11868 45052 11868 45052 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 11132 45052 11132 45052 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 11132 45052 11132 45052 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 11132 45052 11132 45052 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 11132 45052 11132 45052 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 600 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 10396 45052 10396 45052 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 10396 45052 10396 45052 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 10396 45052 10396 45052 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 10396 45052 10396 45052 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 600 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 9660 45052 9660 45052 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 9660 45052 9660 45052 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 9660 45052 9660 45052 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 9660 45052 9660 45052 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 8924 45052 8924 45052 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 8924 45052 8924 45052 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 8924 45052 8924 45052 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 8924 45052 8924 45052 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 600 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 8188 45052 8188 45052 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 8188 45052 8188 45052 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 8188 45052 8188 45052 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 8188 45052 8188 45052 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 600 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 7452 45052 7452 45052 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 7452 45052 7452 45052 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 7452 45052 7452 45052 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 7452 45052 7452 45052 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 6716 45052 6716 45052 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 6716 45052 6716 45052 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 6716 45052 6716 45052 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 6716 45052 6716 45052 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 17756 45052 17756 45052 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 17756 45052 17756 45052 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 17756 45052 17756 45052 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 17756 45052 17756 45052 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 600 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 17020 45052 17020 45052 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 17020 45052 17020 45052 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 17020 45052 17020 45052 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 17020 45052 17020 45052 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 600 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 16284 45052 16284 45052 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 16284 45052 16284 45052 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 16284 45052 16284 45052 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 16284 45052 16284 45052 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 15548 45052 15548 45052 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 15548 45052 15548 45052 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 15548 45052 15548 45052 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 15548 45052 15548 45052 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 600 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 14812 45052 14812 45052 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 14812 45052 14812 45052 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 14812 45052 14812 45052 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 14812 45052 14812 45052 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 600 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 14076 45052 14076 45052 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 14076 45052 14076 45052 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 14076 45052 14076 45052 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 14076 45052 14076 45052 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 13340 45052 13340 45052 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 13340 45052 13340 45052 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 13340 45052 13340 45052 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 13340 45052 13340 45052 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 600 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 12604 45052 12604 45052 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 12604 45052 12604 45052 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 12604 45052 12604 45052 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 12604 45052 12604 45052 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 200 1000 500 44152 1 FreeSans 6000 0 0 0 VPWR
port 52 nsew
flabel metal4 s 9800 1000 10100 44152 1 FreeSans 6000 0 0 0 VGND
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
